<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-57.2314,-59.5427,96.7078,-140.3</PageViewport>
<gate>
<ID>1</ID>
<type>DE_TO</type>
<position>144,-150.5</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R39</lparam></gate>
<gate>
<ID>2</ID>
<type>DA_FROM</type>
<position>99.5,-36.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_AND2</type>
<position>81,84</position>
<input>
<ID>IN_0</ID>102 </input>d
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>104.5,-31.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>144,-161</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R47</lparam></gate>
<gate>
<ID>6</ID>
<type>EE_VDD</type>
<position>107.5,-37</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>80,91</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_MUX_8x1</type>
<position>6.5,-17.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>3 </input>
<input>
<ID>IN_4</ID>25 </input>
<input>
<ID>IN_5</ID>26 </input>
<input>
<ID>IN_6</ID>27 </input>
<input>
<ID>IN_7</ID>28 </input>
<output>
<ID>OUT</ID>130 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>9</ID>
<type>FF_GND</type>
<position>107.5,-34</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AI_MUX_8x1</type>
<position>61,-17.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>84 </input>
<input>
<ID>IN_4</ID>85 </input>
<input>
<ID>IN_5</ID>125 </input>
<input>
<ID>IN_6</ID>87 </input>
<input>
<ID>IN_7</ID>88 </input>
<output>
<ID>OUT</ID>138 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>143.5,-172.5</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R55</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>112.5,-34</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>82,91</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>113,-37</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>-18,54</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_MUX_2x1</type>
<position>78.5,-64.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>378 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_MUX_2x1</type>
<position>84.5,-64.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>379 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AI_MUX_8x1</type>
<position>92.5,-35</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>4 </input>
<input>
<ID>IN_6</ID>4 </input>
<input>
<ID>IN_7</ID>5 </input>
<output>
<ID>OUT</ID>143 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_MUX_2x1</type>
<position>90,-64.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>380 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_FULLADDER_4BIT</type>
<position>53,-42</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>134 </input>
<input>
<ID>IN_3</ID>130 </input>
<input>
<ID>IN_B_0</ID>135 </input>
<input>
<ID>IN_B_1</ID>136 </input>
<input>
<ID>IN_B_2</ID>137 </input>
<input>
<ID>IN_B_3</ID>138 </input>
<output>
<ID>OUT_0</ID>165 </output>
<output>
<ID>OUT_1</ID>164 </output>
<output>
<ID>OUT_2</ID>166 </output>
<output>
<ID>OUT_3</ID>167 </output>
<input>
<ID>carry_in</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_MUX_2x1</type>
<position>95.5,-64.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>381 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>-2,-0.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_MUX_2x1</type>
<position>101,-64.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>382 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>2.5,-2.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_MUX_2x1</type>
<position>106.5,-66</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>383 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>5.5,-4</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_MUX_2x1</type>
<position>112,-64.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>384 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_MUX_2x1</type>
<position>117.5,-64.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>385 </output>
<input>
<ID>SEL_0</ID>8 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>-19,61</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>129.5,-63.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID S3</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>-17,61</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>77.5,-60.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU0</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>79.5,-60.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>83.5,-60.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU1</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>85.5,-60.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>89,-60</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU2</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>91,-60</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>94.5,-60.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU3</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>97,-60.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>100,-60.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>102,-60.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M4</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>105.5,-60.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>-4.5,-12</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-3,6</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>-1,6</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>1.5,4</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>3.5,4</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>5.5,4</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>107.5,-60.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M5</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>111,-60.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>113,-60.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M6</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>116.5,-60.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>119,-60.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M7</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>-13.5,54</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>7,-7.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>8,-12.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>9,-7.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>11.5,-12.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>59</ID>
<type>AI_MUX_8x1</type>
<position>20.5,-17.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_2</ID>30 </input>
<input>
<ID>IN_3</ID>31 </input>
<input>
<ID>IN_4</ID>38 </input>
<input>
<ID>IN_5</ID>39 </input>
<input>
<ID>IN_6</ID>40 </input>
<input>
<ID>IN_7</ID>41 </input>
<output>
<ID>OUT</ID>134 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>12,-0.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_OR2</type>
<position>16.5,-2.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_SMALL_INVERTER</type>
<position>20,-3</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>14,-11.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>11,5.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>13,6.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>15.5,5.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>17.5,3.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>20.5,4.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>21,-7.5</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>22,-12.5</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>23,-7.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>24,-12.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>73</ID>
<type>AI_MUX_8x1</type>
<position>34,-18.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>43 </input>
<input>
<ID>IN_3</ID>44 </input>
<input>
<ID>IN_4</ID>51 </input>
<input>
<ID>IN_5</ID>52 </input>
<input>
<ID>IN_6</ID>53 </input>
<input>
<ID>IN_7</ID>54 </input>
<output>
<ID>OUT</ID>133 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>25.5,-1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_OR2</type>
<position>30,-3</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_SMALL_INVERTER</type>
<position>33.5,-3.5</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>27.5,-12</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>24.5,6.5</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>26.5,6</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>29,4</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>31,3</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>33.5,1</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>34.5,-8</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>35.5,-13</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>36.5,-8</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>37.5,-13</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>87</ID>
<type>AI_MUX_8x1</type>
<position>48,-18</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>56 </input>
<input>
<ID>IN_3</ID>57 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>66 </input>
<input>
<ID>IN_7</ID>67 </input>
<output>
<ID>OUT</ID>132 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>39.5,-1</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_OR2</type>
<position>44,-3</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_SMALL_INVERTER</type>
<position>47.5,-3</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>41.5,-12</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>38.5,5.5</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>40.5,5</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>43,2.5</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>45,3</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>47.5,1.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>48.5,-8.5</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>50.5,-10.5</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>52,-4.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>53.5,-11.5</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>-14.5,61</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>56,-5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>-12.5,61</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND2</type>
<position>-9,54</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>-10,61</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_FULLADDER_4BIT</type>
<position>3,40</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_2</ID>192 </input>
<input>
<ID>IN_3</ID>193 </input>
<input>
<ID>IN_B_0</ID>237 </input>
<input>
<ID>IN_B_1</ID>236 </input>
<input>
<ID>IN_B_2</ID>235 </input>
<input>
<ID>IN_B_3</ID>234 </input>
<output>
<ID>OUT_0</ID>239 </output>
<output>
<ID>OUT_1</ID>240 </output>
<output>
<ID>OUT_2</ID>241 </output>
<output>
<ID>OUT_3</ID>242 </output>
<input>
<ID>carry_in</ID>238 </input>
<output>
<ID>carry_out</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>107</ID>
<type>DA_FROM</type>
<position>-8,61</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>144,-184</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R63</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>-4,54</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>175,-103</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R8</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>-5,61</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>-3,61</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>174.5,-114</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>173.5,-125</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R24</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>174,-135</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R32</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>174,-150</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R40</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>174,-161</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R48</lparam></gate>
<gate>
<ID>118</ID>
<type>DA_FROM</type>
<position>58,-9.5</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>59.5,-5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>60.5,-11</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>61.5,-7</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>62.5,7.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>63.5,-8</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>64.5,-12</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>125</ID>
<type>AI_MUX_8x1</type>
<position>74.5,-17</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_4</ID>93 </input>
<input>
<ID>IN_5</ID>126 </input>
<input>
<ID>IN_6</ID>95 </input>
<input>
<ID>IN_7</ID>96 </input>
<output>
<ID>OUT</ID>137 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>69.5,-4.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>71.5,-9</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>72.5,-4.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>74,-10.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>75,-6.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>76,8</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>77,-7.5</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>78,-11.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AI_MUX_8x1</type>
<position>87,-16.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>99 </input>
<input>
<ID>IN_3</ID>100 </input>
<input>
<ID>IN_4</ID>101 </input>
<input>
<ID>IN_5</ID>127 </input>
<input>
<ID>IN_6</ID>129 </input>
<input>
<ID>IN_7</ID>104 </input>
<output>
<ID>OUT</ID>136 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>82,-4</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>84,-8.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>85.5,-4</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>86.5,-10</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>87.5,-6</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>173.5,-171.5</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R56</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>89,8.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>93,-9.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>143</ID>
<type>AI_MUX_8x1</type>
<position>101,-16.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>107 </input>
<input>
<ID>IN_3</ID>108 </input>
<input>
<ID>IN_4</ID>109 </input>
<input>
<ID>IN_5</ID>128 </input>
<input>
<ID>IN_6</ID>111 </input>
<input>
<ID>IN_7</ID>112 </input>
<output>
<ID>OUT</ID>135 </output>
<input>
<ID>SEL_0</ID>142 </input>
<input>
<ID>SEL_1</ID>141 </input>
<input>
<ID>SEL_2</ID>139 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>96,-4</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>98,-8.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>99.5,-4</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>100.5,-10</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>101.5,-6</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>102.5,8</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>103.5,-7</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>106.5,-8</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 1</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>173.5,-182</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R64</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_DFF_LOW</type>
<position>-28,-108.5</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>315 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>119 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>-37,-109.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_DFF_LOW</type>
<position>-27.5,-119</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>316 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>120 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>-37.5,-118.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_DFF_LOW</type>
<position>-28,-130</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>317 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>131 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>-37.5,-130.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>159</ID>
<type>AE_DFF_LOW</type>
<position>-28,-140.5</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>318 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>273 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>-35,-141.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_DFF_LOW</type>
<position>-2.5,-108</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>322 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>140 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_SMALL_INVERTER</type>
<position>62.5,2</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>76,3</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>89,3.5</position>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>102.5,2.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>-9,-110</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_DFF_LOW</type>
<position>-2.5,-119</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>323 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>168 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>DA_FROM</type>
<position>-9,-120.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>90,-7</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_DFF_LOW</type>
<position>-3,-130</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>324 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>169 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>-4.5,-24.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>-10,-26.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>-4.5,-31</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>-11.5,-131.5</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>175</ID>
<type>DD_KEYPAD_HEX</type>
<position>-17.5,-50.5</position>
<output>
<ID>OUT_0</ID>147 </output>
<output>
<ID>OUT_1</ID>146 </output>
<output>
<ID>OUT_2</ID>145 </output>
<output>
<ID>OUT_3</ID>144 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_DFF_LOW</type>
<position>-3,-140.5</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>325 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>280 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>-11,-142</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-107.5</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>330 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>170 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>14.5,-108.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_DFF_LOW</type>
<position>24,-118</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>331 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>171 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>181</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>174.5,-70.5</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>392 </input>
<input>
<ID>IN_2</ID>391 </input>
<input>
<ID>IN_3</ID>390 </input>
<input>
<ID>IN_4</ID>389 </input>
<input>
<ID>IN_5</ID>388 </input>
<input>
<ID>IN_6</ID>387 </input>
<input>
<ID>IN_7</ID>386 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>18,-119</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-129</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>332 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>172 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>15,-130.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>185</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>31.5,-71.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>157 </input>
<input>
<ID>IN_3</ID>156 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-139.5</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>333 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>281 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>-5.5,-44</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S3</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>-6.5,-49</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>-4.5,-52</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>-7,-55.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>191</ID>
<type>DD_KEYPAD_HEX</type>
<position>6,-50</position>
<output>
<ID>OUT_0</ID>151 </output>
<output>
<ID>OUT_1</ID>150 </output>
<output>
<ID>OUT_2</ID>149 </output>
<output>
<ID>OUT_3</ID>148 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>192</ID>
<type>DE_TO</type>
<position>17,-44</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>193</ID>
<type>DE_TO</type>
<position>16,-49</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>194</ID>
<type>DE_TO</type>
<position>18,-51.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>195</ID>
<type>DE_TO</type>
<position>15.5,-55.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>196</ID>
<type>DD_KEYPAD_HEX</type>
<position>25,-50</position>
<output>
<ID>OUT_0</ID>155 </output>
<output>
<ID>OUT_1</ID>154 </output>
<output>
<ID>OUT_2</ID>153 </output>
<output>
<ID>OUT_3</ID>152 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>197</ID>
<type>DE_TO</type>
<position>37.5,-44</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>198</ID>
<type>DE_TO</type>
<position>36.5,-49</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>38.5,-51.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>200</ID>
<type>DE_TO</type>
<position>36,-55.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>16.5,-140.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>19,-67</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>19.5,-70</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>16.5,-71.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>17.5,-74.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>45.5,-66</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>46,-69</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>43,-70.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>44,-73.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>210</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>58,-70.5</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>161 </input>
<input>
<ID>IN_3</ID>160 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-106.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>338 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>173 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>53,-51.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU1</lparam></gate>
<gate>
<ID>213</ID>
<type>DE_TO</type>
<position>55.5,-52.5</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU0</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>50.5,-54</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU2</lparam></gate>
<gate>
<ID>215</ID>
<type>DE_TO</type>
<position>46.5,-52.5</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ALU3</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>46.5,-108</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_DFF_LOW</type>
<position>53,-117</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>339 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>174 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>45,-118</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-128</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>340 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>175 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>7,74</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>DA_FROM</type>
<position>6,81</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>8,81</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND2</type>
<position>11.5,74</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>10.5,81</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>12.5,81</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_AND2</type>
<position>16,74</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>15,81</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_FULLADDER_4BIT</type>
<position>28,60</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<input>
<ID>IN_2</ID>204 </input>
<input>
<ID>IN_3</ID>205 </input>
<input>
<ID>IN_B_0</ID>248 </input>
<input>
<ID>IN_B_1</ID>247 </input>
<input>
<ID>IN_B_2</ID>246 </input>
<input>
<ID>IN_B_3</ID>245 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>237 </output>
<output>
<ID>OUT_2</ID>236 </output>
<output>
<ID>OUT_3</ID>235 </output>
<input>
<ID>carry_in</ID>253 </input>
<output>
<ID>carry_out</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>17,81</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>21,74</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>20,81</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>22,81</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>35,85.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>34,92.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>36,92.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>39.5,85.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>38.5,92.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>40.5,92.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>44,85.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>43,92.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_FULLADDER_4BIT</type>
<position>56,71.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>215 </input>
<input>
<ID>IN_2</ID>216 </input>
<input>
<ID>IN_3</ID>217 </input>
<input>
<ID>IN_B_0</ID>230 </input>
<input>
<ID>IN_B_1</ID>232 </input>
<input>
<ID>IN_B_2</ID>231 </input>
<input>
<ID>IN_B_3</ID>252 </input>
<output>
<ID>OUT_0</ID>249 </output>
<output>
<ID>OUT_1</ID>248 </output>
<output>
<ID>OUT_2</ID>247 </output>
<output>
<ID>OUT_3</ID>246 </output>
<input>
<ID>carry_in</ID>250 </input>
<output>
<ID>carry_out</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>45,92.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>49,85.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>48,92.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>50,92.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>46.5,-128.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>247</ID>
<type>AE_DFF_LOW</type>
<position>52,-138.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>341 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>282 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>43.5,-140</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_AND2</type>
<position>63,89.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>62,96.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>64,96.5</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_AND2</type>
<position>67.5,89.5</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>66.5,96.5</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_DFF_LOW</type>
<position>84,-105.5</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>346 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>176 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>68.5,96.5</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>72.5,89.5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>71.5,96.5</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>73.5,96.5</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>76,-107</position>
<input>
<ID>IN_0</ID>176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>14,41</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>261</ID>
<type>AE_DFF_LOW</type>
<position>84.5,-116</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>347 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>177 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>262</ID>
<type>DE_TO</type>
<position>6,28</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<gate>
<ID>263</ID>
<type>DA_FROM</type>
<position>76.5,-117</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>264</ID>
<type>DE_TO</type>
<position>3.5,28</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M4</lparam></gate>
<gate>
<ID>265</ID>
<type>AE_DFF_LOW</type>
<position>84,-127</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>348 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>178 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>266</ID>
<type>DE_TO</type>
<position>2,23</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M5</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>77.5,-128</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>268</ID>
<type>DE_TO</type>
<position>-1,25</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M6</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_DFF_LOW</type>
<position>84,-137.5</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>349 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>283 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>270</ID>
<type>DE_TO</type>
<position>-6,26</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M7</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>73,-139</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>272</ID>
<type>DE_TO</type>
<position>30,48.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>273</ID>
<type>AE_DFF_LOW</type>
<position>111,-105</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>354 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>179 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>57.5,63.5</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>275</ID>
<type>DA_FROM</type>
<position>106,-106</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>276</ID>
<type>DA_FROM</type>
<position>66,72.5</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>277</ID>
<type>AE_DFF_LOW</type>
<position>111.5,-115.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>355 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>180 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>278</ID>
<type>DE_TO</type>
<position>81,78.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>279</ID>
<type>DA_FROM</type>
<position>106,-116.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>280</ID>
<type>DA_FROM</type>
<position>58,84.5</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>281</ID>
<type>AE_DFF_LOW</type>
<position>111,-126.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>356 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>181 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>40,60.5</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>103,-127.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>284</ID>
<type>AE_DFF_LOW</type>
<position>111,-137</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>357 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>284 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>102.5,-138.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_DFF_LOW</type>
<position>137.5,-104.5</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>362 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>182 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>132,-105</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_DFF_LOW</type>
<position>138,-115</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>363 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>183 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>130.5,-115</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_DFF_LOW</type>
<position>137.5,-126</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>364 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>184 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>130.5,-126.5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_DFF_LOW</type>
<position>137.5,-136.5</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>365 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>285 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>293</ID>
<type>DA_FROM</type>
<position>130,-137</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_DFF_LOW</type>
<position>165.5,-105.5</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>370 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>185 </input>
<input>
<ID>set</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>158.5,-106.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>296</ID>
<type>AE_DFF_LOW</type>
<position>165.5,-116</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>371 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>186 </input>
<input>
<ID>set</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>159,-115.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>298</ID>
<type>AE_DFF_LOW</type>
<position>166,-127</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>372 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>187 </input>
<input>
<ID>set</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>159,-126.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_DFF_LOW</type>
<position>165.5,-137</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>373 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>270 </input>
<input>
<ID>set</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>301</ID>
<type>DA_FROM</type>
<position>158.5,-137.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_DFF_LOW</type>
<position>164.5,-152</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>374 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>188 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>157,-153</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_DFF_LOW</type>
<position>165,-162.5</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>375 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>189 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>159.5,-163.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>164.5,-173.5</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>376 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>218 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>157.5,-174</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_DFF_LOW</type>
<position>164.5,-184</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>377 </output>
<input>
<ID>clear</ID>314 </input>
<input>
<ID>clock</ID>271 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>157,-185.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>310</ID>
<type>AE_DFF_LOW</type>
<position>137,-152</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>366 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>219 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>129.5,-153</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_DFF_LOW</type>
<position>137.5,-162.5</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>367 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>226 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>130,-163.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_DFF_LOW</type>
<position>137,-173.5</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>368 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>227 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>130,-174.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>316</ID>
<type>AE_DFF_LOW</type>
<position>137,-184</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>369 </output>
<input>
<ID>clear</ID>313 </input>
<input>
<ID>clock</ID>272 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>128.5,-184</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_DFF_LOW</type>
<position>111,-151.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>358 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>228 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>102.5,-154</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_DFF_LOW</type>
<position>111.5,-162</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>359 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>229 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>104.5,-163</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_DFF_LOW</type>
<position>111,-173</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>360 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>233 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>103,-174</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_DFF_LOW</type>
<position>111,-183.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>361 </output>
<input>
<ID>clear</ID>312 </input>
<input>
<ID>clock</ID>279 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>DA_FROM</type>
<position>103.5,-185</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_DFF_LOW</type>
<position>83,-152</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>350 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>254 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>76,-153</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_DFF_LOW</type>
<position>83.5,-162.5</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>351 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>255 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>71.5,-164.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>330</ID>
<type>AE_DFF_LOW</type>
<position>82.5,-173.5</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>352 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>256 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>72.5,-174.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_DFF_LOW</type>
<position>82.5,-184</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>353 </output>
<input>
<ID>clear</ID>311 </input>
<input>
<ID>clock</ID>278 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>75.5,-185.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_DFF_LOW</type>
<position>24,-154</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>334 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>257 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>335</ID>
<type>DA_FROM</type>
<position>15.5,-154</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>24.5,-164</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>335 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>258 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>16.5,-164</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_DFF_LOW</type>
<position>24,-175</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>336 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>259 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>339</ID>
<type>DA_FROM</type>
<position>18.5,-176</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>340</ID>
<type>AE_DFF_LOW</type>
<position>24,-185.5</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>337 </output>
<input>
<ID>clear</ID>309 </input>
<input>
<ID>clock</ID>276 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>14.5,-186.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-152.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>342 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>260 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>44,-153.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_DFF_LOW</type>
<position>53,-163</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>343 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>261 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>45,-164</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-174</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>344 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>262 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>45.5,-175.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>348</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-184.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>345 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>277 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>45.5,-185</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_DFF_LOW</type>
<position>-3,-153</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>326 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>263 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>-8.5,-154</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>352</ID>
<type>AE_DFF_LOW</type>
<position>-2.5,-163.5</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>327 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>264 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>-9.5,-164.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>354</ID>
<type>AE_DFF_LOW</type>
<position>-3,-174.5</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>328 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>265 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>355</ID>
<type>DA_FROM</type>
<position>-9.5,-175</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_DFF_LOW</type>
<position>-3,-185</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>329 </output>
<input>
<ID>clear</ID>308 </input>
<input>
<ID>clock</ID>275 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>-14.5,-185.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_DFF_LOW</type>
<position>-28,-153</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>319 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>266 </input>
<input>
<ID>set</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>-34.5,-154.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_DFF_LOW</type>
<position>-27.5,-163.5</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>320 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>267 </input>
<input>
<ID>set</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>-34.5,-164.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>362</ID>
<type>AE_DFF_LOW</type>
<position>-28,-174.5</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>321 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>268 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>363</ID>
<type>DA_FROM</type>
<position>-36,-175.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_DFF_LOW</type>
<position>-28,-185</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>307 </output>
<input>
<ID>clear</ID>307 </input>
<input>
<ID>clock</ID>274 </input>
<input>
<ID>set</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>365</ID>
<type>DA_FROM</type>
<position>-36,-184.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>366</ID>
<type>BE_DECODER_3x8</type>
<position>-65,-132.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>306 </input>
<input>
<ID>IN_2</ID>304 </input>
<output>
<ID>OUT_0</ID>292 </output>
<output>
<ID>OUT_1</ID>291 </output>
<output>
<ID>OUT_2</ID>290 </output>
<output>
<ID>OUT_3</ID>289 </output>
<output>
<ID>OUT_4</ID>288 </output>
<output>
<ID>OUT_5</ID>287 </output>
<output>
<ID>OUT_6</ID>286 </output>
<output>
<ID>OUT_7</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>368</ID>
<type>AA_RAM_4x4</type>
<position>-84.5,-166.5</position>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_TOGGLE</type>
<position>-54.5,-66</position>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>376</ID>
<type>BB_CLOCK</type>
<position>-56,-72.5</position>
<output>
<ID>CLK</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>377</ID>
<type>DE_TO</type>
<position>-50,-72.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clock</lparam></gate>
<gate>
<ID>378</ID>
<type>DE_TO</type>
<position>-47.5,-66</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_TOGGLE</type>
<position>-72.5,-132.5</position>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_TOGGLE</type>
<position>-73,-139.5</position>
<output>
<ID>OUT_0</ID>305 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_TOGGLE</type>
<position>-76,-135</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>383</ID>
<type>DA_FROM</type>
<position>-24.5,-197</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>5,-197</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>28.5,-194.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>60,-195</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>87.5,-195</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>116,-194</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>144,-194.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>175.5,-195</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O</lparam></gate>
<gate>
<ID>391</ID>
<type>DE_TO</type>
<position>-21,-106</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1</lparam></gate>
<gate>
<ID>392</ID>
<type>DE_TO</type>
<position>-18,-117.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R9</lparam></gate>
<gate>
<ID>393</ID>
<type>DE_TO</type>
<position>-19,-128</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17</lparam></gate>
<gate>
<ID>394</ID>
<type>DE_TO</type>
<position>-19,-139.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R25</lparam></gate>
<gate>
<ID>395</ID>
<type>DE_TO</type>
<position>-19,-151</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R33</lparam></gate>
<gate>
<ID>396</ID>
<type>DE_TO</type>
<position>-19.5,-162.5</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R41</lparam></gate>
<gate>
<ID>397</ID>
<type>DE_TO</type>
<position>-19,-173</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R49</lparam></gate>
<gate>
<ID>398</ID>
<type>DE_TO</type>
<position>-17.5,-183</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R57</lparam></gate>
<gate>
<ID>399</ID>
<type>DE_TO</type>
<position>5.5,-106</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R2</lparam></gate>
<gate>
<ID>400</ID>
<type>DE_TO</type>
<position>4,-117</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R10</lparam></gate>
<gate>
<ID>401</ID>
<type>DE_TO</type>
<position>3.5,-128.5</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R18</lparam></gate>
<gate>
<ID>402</ID>
<type>DE_TO</type>
<position>4.5,-138.5</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R26</lparam></gate>
<gate>
<ID>403</ID>
<type>DE_TO</type>
<position>4,-150.5</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R34</lparam></gate>
<gate>
<ID>404</ID>
<type>DE_TO</type>
<position>4,-161.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R42</lparam></gate>
<gate>
<ID>405</ID>
<type>DE_TO</type>
<position>3.5,-173</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R50</lparam></gate>
<gate>
<ID>406</ID>
<type>DE_TO</type>
<position>3.5,-183.5</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R58</lparam></gate>
<gate>
<ID>407</ID>
<type>DE_TO</type>
<position>31,-104.5</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R3</lparam></gate>
<gate>
<ID>408</ID>
<type>DE_TO</type>
<position>30.5,-116</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R11</lparam></gate>
<gate>
<ID>409</ID>
<type>DE_TO</type>
<position>31,-126</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R19</lparam></gate>
<gate>
<ID>410</ID>
<type>DE_TO</type>
<position>31,-137</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R27</lparam></gate>
<gate>
<ID>411</ID>
<type>DE_TO</type>
<position>31,-151.5</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R35</lparam></gate>
<gate>
<ID>412</ID>
<type>DE_TO</type>
<position>31.5,-162</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R43</lparam></gate>
<gate>
<ID>413</ID>
<type>DE_TO</type>
<position>31.5,-172.5</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R51</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_TO</type>
<position>32,-183.5</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R59</lparam></gate>
<gate>
<ID>415</ID>
<type>DE_TO</type>
<position>61,-105</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R4</lparam></gate>
<gate>
<ID>416</ID>
<type>DE_TO</type>
<position>60,-115</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R12</lparam></gate>
<gate>
<ID>417</ID>
<type>DE_TO</type>
<position>60.5,-126</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R20</lparam></gate>
<gate>
<ID>418</ID>
<type>DE_TO</type>
<position>60,-136.5</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R28</lparam></gate>
<gate>
<ID>419</ID>
<type>DE_TO</type>
<position>59.5,-151</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R36</lparam></gate>
<gate>
<ID>420</ID>
<type>DE_TO</type>
<position>60,-160.5</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R44</lparam></gate>
<gate>
<ID>421</ID>
<type>DE_TO</type>
<position>60,-171.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R52</lparam></gate>
<gate>
<ID>422</ID>
<type>DE_TO</type>
<position>59.5,-181.5</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R60</lparam></gate>
<gate>
<ID>423</ID>
<type>DE_TO</type>
<position>91,-105</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R5</lparam></gate>
<gate>
<ID>424</ID>
<type>DE_TO</type>
<position>92,-114</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R13</lparam></gate>
<gate>
<ID>425</ID>
<type>DE_TO</type>
<position>92.5,-124.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R21</lparam></gate>
<gate>
<ID>426</ID>
<type>DE_TO</type>
<position>91.5,-135.5</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R29</lparam></gate>
<gate>
<ID>427</ID>
<type>DE_TO</type>
<position>91.5,-149.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R37</lparam></gate>
<gate>
<ID>428</ID>
<type>DE_TO</type>
<position>90.5,-160</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R45</lparam></gate>
<gate>
<ID>429</ID>
<type>DE_TO</type>
<position>91,-171</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R53</lparam></gate>
<gate>
<ID>430</ID>
<type>DE_TO</type>
<position>90.5,-181.5</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R61</lparam></gate>
<gate>
<ID>431</ID>
<type>DE_TO</type>
<position>118,-103.5</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R6</lparam></gate>
<gate>
<ID>432</ID>
<type>DE_TO</type>
<position>118.5,-113.5</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R14</lparam></gate>
<gate>
<ID>433</ID>
<type>DE_TO</type>
<position>117,-125</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R22</lparam></gate>
<gate>
<ID>434</ID>
<type>DE_TO</type>
<position>118.5,-137</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R30</lparam></gate>
<gate>
<ID>435</ID>
<type>DE_TO</type>
<position>118.5,-149</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R38</lparam></gate>
<gate>
<ID>436</ID>
<type>DE_TO</type>
<position>117.5,-160</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R46</lparam></gate>
<gate>
<ID>437</ID>
<type>DE_TO</type>
<position>118,-171.5</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R54</lparam></gate>
<gate>
<ID>438</ID>
<type>DE_TO</type>
<position>118,-181</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R62</lparam></gate>
<gate>
<ID>439</ID>
<type>DE_TO</type>
<position>143.5,-104</position>
<input>
<ID>IN_0</ID>362 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R7</lparam></gate>
<gate>
<ID>440</ID>
<type>DE_TO</type>
<position>145,-113.5</position>
<input>
<ID>IN_0</ID>363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R15</lparam></gate>
<gate>
<ID>441</ID>
<type>DE_TO</type>
<position>144.5,-124.5</position>
<input>
<ID>IN_0</ID>364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R23</lparam></gate>
<gate>
<ID>442</ID>
<type>DE_TO</type>
<position>144.5,-135</position>
<input>
<ID>IN_0</ID>365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R31</lparam></gate>
<gate>
<ID>444</ID>
<type>DE_TO</type>
<position>78.5,-73.5</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT1</lparam></gate>
<gate>
<ID>445</ID>
<type>DE_TO</type>
<position>84.5,-73.5</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT2</lparam></gate>
<gate>
<ID>446</ID>
<type>DE_TO</type>
<position>90,-74</position>
<input>
<ID>IN_0</ID>380 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT3</lparam></gate>
<gate>
<ID>447</ID>
<type>DE_TO</type>
<position>95.5,-73.5</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT4</lparam></gate>
<gate>
<ID>448</ID>
<type>DE_TO</type>
<position>101,-73.5</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT5</lparam></gate>
<gate>
<ID>449</ID>
<type>DE_TO</type>
<position>106.5,-74</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT6</lparam></gate>
<gate>
<ID>450</ID>
<type>DE_TO</type>
<position>112,-74</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT7</lparam></gate>
<gate>
<ID>451</ID>
<type>DE_TO</type>
<position>117.5,-73.5</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT8</lparam></gate>
<gate>
<ID>453</ID>
<type>DA_FROM</type>
<position>156.5,-66</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT8</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>158,-68.5</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT7</lparam></gate>
<gate>
<ID>455</ID>
<type>DA_FROM</type>
<position>156,-71</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT6</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>155,-75</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT5</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>154.5,-79</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT4</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>158,-82</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT3</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>163,-85</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPUT2</lparam></gate>
<gate>
<ID>460</ID>
<type>DA_FROM</type>
<position>168.5,-82</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID INPUT1</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>-33.5,-89.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT1</lparam></gate>
<gate>
<ID>463</ID>
<type>DA_FROM</type>
<position>-11.5,-87.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT2</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>14.5,-87.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT3</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>40,-89</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT4</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>70.5,-88.5</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT5</lparam></gate>
<gate>
<ID>467</ID>
<type>DA_FROM</type>
<position>101.5,-92</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT6</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>127.5,-90</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT7</lparam></gate>
<gate>
<ID>469</ID>
<type>DA_FROM</type>
<position>146.5,-91.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID INPUT8</lparam></gate>
<gate>
<ID>471</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>118,-208</position>
<input>
<ID>IN_0</ID>401 </input>
<input>
<ID>IN_1</ID>400 </input>
<input>
<ID>IN_2</ID>399 </input>
<input>
<ID>IN_3</ID>398 </input>
<input>
<ID>IN_4</ID>397 </input>
<input>
<ID>IN_5</ID>396 </input>
<input>
<ID>IN_6</ID>395 </input>
<input>
<ID>IN_7</ID>394 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>108.5,-202</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R8</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>106,-205</position>
<input>
<ID>IN_0</ID>395 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R7</lparam></gate>
<gate>
<ID>475</ID>
<type>DA_FROM</type>
<position>94.5,-205.5</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R6</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>91.5,-207.5</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R5</lparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>98,-208.5</position>
<input>
<ID>IN_0</ID>398 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R4</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>106.5,-210</position>
<input>
<ID>IN_0</ID>399 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R3</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>107,-213</position>
<input>
<ID>IN_0</ID>400 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R2</lparam></gate>
<gate>
<ID>480</ID>
<type>DA_FROM</type>
<position>108.5,-216</position>
<input>
<ID>IN_0</ID>401 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1</lparam></gate>
<gate>
<ID>482</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>118.5,-228</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>408 </input>
<input>
<ID>IN_2</ID>407 </input>
<input>
<ID>IN_3</ID>406 </input>
<input>
<ID>IN_4</ID>405 </input>
<input>
<ID>IN_5</ID>404 </input>
<input>
<ID>IN_6</ID>403 </input>
<input>
<ID>IN_7</ID>402 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>483</ID>
<type>DA_FROM</type>
<position>107.5,-222</position>
<input>
<ID>IN_0</ID>402 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16</lparam></gate>
<gate>
<ID>484</ID>
<type>DA_FROM</type>
<position>103,-224.5</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R15</lparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>100,-226</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R14</lparam></gate>
<gate>
<ID>486</ID>
<type>DA_FROM</type>
<position>106.5,-227.5</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R13</lparam></gate>
<gate>
<ID>487</ID>
<type>DA_FROM</type>
<position>96.5,-229</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R12</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>107,-230</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R11</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>107.5,-233</position>
<input>
<ID>IN_0</ID>408 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R10</lparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>112,-236</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R9</lparam></gate>
<gate>
<ID>491</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>119,-246</position>
<input>
<ID>IN_0</ID>417 </input>
<input>
<ID>IN_1</ID>416 </input>
<input>
<ID>IN_2</ID>415 </input>
<input>
<ID>IN_3</ID>414 </input>
<input>
<ID>IN_4</ID>413 </input>
<input>
<ID>IN_5</ID>412 </input>
<input>
<ID>IN_6</ID>411 </input>
<input>
<ID>IN_7</ID>410 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>111,-242</position>
<input>
<ID>IN_0</ID>410 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R24</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>104,-243.5</position>
<input>
<ID>IN_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R23</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>95.5,-243</position>
<input>
<ID>IN_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R22</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>107,-245.5</position>
<input>
<ID>IN_0</ID>413 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R21</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>99,-246.5</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R20</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>102.5,-248.5</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R19</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>108,-251</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R18</lparam></gate>
<gate>
<ID>499</ID>
<type>DA_FROM</type>
<position>112.5,-254</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17</lparam></gate>
<gate>
<ID>500</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>119,-262.5</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>424 </input>
<input>
<ID>IN_2</ID>423 </input>
<input>
<ID>IN_3</ID>422 </input>
<input>
<ID>IN_4</ID>421 </input>
<input>
<ID>IN_5</ID>420 </input>
<input>
<ID>IN_6</ID>419 </input>
<input>
<ID>IN_7</ID>418 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>501</ID>
<type>DA_FROM</type>
<position>111,-258.5</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R32</lparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>107,-259.5</position>
<input>
<ID>IN_0</ID>419 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R31</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>100.5,-260.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R30</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>107,-262</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R29</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>99.5,-263.5</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R28</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>107.5,-264.5</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R27</lparam></gate>
<gate>
<ID>507</ID>
<type>DA_FROM</type>
<position>108,-267.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R26</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>112.5,-270.5</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R25</lparam></gate>
<gate>
<ID>509</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>119.5,-281</position>
<input>
<ID>IN_0</ID>433 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>431 </input>
<input>
<ID>IN_3</ID>430 </input>
<input>
<ID>IN_4</ID>429 </input>
<input>
<ID>IN_5</ID>428 </input>
<input>
<ID>IN_6</ID>427 </input>
<input>
<ID>IN_7</ID>426 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>110.5,-275.5</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R40</lparam></gate>
<gate>
<ID>511</ID>
<type>DA_FROM</type>
<position>107.5,-278</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R39</lparam></gate>
<gate>
<ID>512</ID>
<type>DA_FROM</type>
<position>101,-279</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R38</lparam></gate>
<gate>
<ID>513</ID>
<type>DA_FROM</type>
<position>107.5,-280.5</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R37</lparam></gate>
<gate>
<ID>514</ID>
<type>DA_FROM</type>
<position>100.5,-281</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R36</lparam></gate>
<gate>
<ID>515</ID>
<type>DA_FROM</type>
<position>108,-283</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R35</lparam></gate>
<gate>
<ID>516</ID>
<type>DA_FROM</type>
<position>108.5,-286</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R34</lparam></gate>
<gate>
<ID>517</ID>
<type>DA_FROM</type>
<position>113,-289</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R33</lparam></gate>
<gate>
<ID>518</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>119.5,-300.5</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>440 </input>
<input>
<ID>IN_2</ID>439 </input>
<input>
<ID>IN_3</ID>438 </input>
<input>
<ID>IN_4</ID>437 </input>
<input>
<ID>IN_5</ID>436 </input>
<input>
<ID>IN_6</ID>435 </input>
<input>
<ID>IN_7</ID>434 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>519</ID>
<type>DA_FROM</type>
<position>111.5,-296.5</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R48</lparam></gate>
<gate>
<ID>520</ID>
<type>DA_FROM</type>
<position>107.5,-297.5</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R47</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>97.5,-298</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R46</lparam></gate>
<gate>
<ID>522</ID>
<type>DA_FROM</type>
<position>107.5,-300</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R45</lparam></gate>
<gate>
<ID>523</ID>
<type>DA_FROM</type>
<position>97.5,-301</position>
<input>
<ID>IN_0</ID>438 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R44</lparam></gate>
<gate>
<ID>524</ID>
<type>DA_FROM</type>
<position>108,-302.5</position>
<input>
<ID>IN_0</ID>439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R43</lparam></gate>
<gate>
<ID>525</ID>
<type>DA_FROM</type>
<position>108.5,-305.5</position>
<input>
<ID>IN_0</ID>440 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R42</lparam></gate>
<gate>
<ID>526</ID>
<type>DA_FROM</type>
<position>113,-308.5</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R41</lparam></gate>
<gate>
<ID>527</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>119.5,-320.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>448 </input>
<input>
<ID>IN_2</ID>447 </input>
<input>
<ID>IN_3</ID>446 </input>
<input>
<ID>IN_4</ID>445 </input>
<input>
<ID>IN_5</ID>444 </input>
<input>
<ID>IN_6</ID>443 </input>
<input>
<ID>IN_7</ID>442 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>528</ID>
<type>DA_FROM</type>
<position>111.5,-315.5</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R56</lparam></gate>
<gate>
<ID>529</ID>
<type>DA_FROM</type>
<position>107.5,-317.5</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R55</lparam></gate>
<gate>
<ID>530</ID>
<type>DA_FROM</type>
<position>101,-318.5</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R54</lparam></gate>
<gate>
<ID>531</ID>
<type>DA_FROM</type>
<position>107.5,-320</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R53</lparam></gate>
<gate>
<ID>532</ID>
<type>DA_FROM</type>
<position>96.5,-320.5</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R52</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>108,-322.5</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R51</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>108.5,-325.5</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R50</lparam></gate>
<gate>
<ID>535</ID>
<type>DA_FROM</type>
<position>113,-328.5</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R49</lparam></gate>
<gate>
<ID>536</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>120.5,-339</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>456 </input>
<input>
<ID>IN_2</ID>455 </input>
<input>
<ID>IN_3</ID>454 </input>
<input>
<ID>IN_4</ID>453 </input>
<input>
<ID>IN_5</ID>452 </input>
<input>
<ID>IN_6</ID>451 </input>
<input>
<ID>IN_7</ID>450 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>112.5,-335</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R64</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>103.5,-334.5</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R63</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>102,-337</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R62</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>108.5,-338.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R61</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>95,-339.5</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R60</lparam></gate>
<gate>
<ID>542</ID>
<type>DA_FROM</type>
<position>109,-341</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R59</lparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>109.5,-344</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R58</lparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>114,-347</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R57</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-9,-2,-3.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3.5,-14.5,3.5,-9</points>
<intersection>-14.5 3</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2,-9,3.5,-9</points>
<intersection>-2 0</intersection>
<intersection>3.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>3.5,-14.5,4,-14.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>3.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-8,2.5,-5.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5,-14.5,5,-8</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-8,5,-8</points>
<intersection>2.5 0</intersection>
<intersection>5 1</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-14.5,5.5,-6</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-14.5,6,-14.5</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-36.5,97.5,-36.5</points>
<connection>
<GID>18</GID>
<name>IN_5</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>97 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>97,-37.5,97,-36.5</points>
<intersection>-37.5 5</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>95.5,-37.5,97,-37.5</points>
<connection>
<GID>18</GID>
<name>IN_6</name></connection>
<intersection>97 4</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-31.5,102.5,-31.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>102 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102,-38.5,102,-31.5</points>
<intersection>-38.5 8</intersection>
<intersection>-35.5 7</intersection>
<intersection>-34.5 6</intersection>
<intersection>-33.5 5</intersection>
<intersection>-32.5 4</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95.5,-32.5,102,-32.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>102 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>95.5,-33.5,102,-33.5</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>102 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>95.5,-34.5,102,-34.5</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<intersection>102 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>95.5,-35.5,102,-35.5</points>
<connection>
<GID>18</GID>
<name>IN_4</name></connection>
<intersection>102 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>95.5,-38.5,102,-38.5</points>
<connection>
<GID>18</GID>
<name>IN_7</name></connection>
<intersection>102 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>108.5,-34,110.5,-34</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-37,111,-37</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-63.5,127.5,-63.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>81 3</intersection>
<intersection>87 4</intersection>
<intersection>92.5 5</intersection>
<intersection>98 6</intersection>
<intersection>103.5 7</intersection>
<intersection>109 8</intersection>
<intersection>114.5 9</intersection>
<intersection>120 10</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-64.5,81,-63.5</points>
<connection>
<GID>16</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>87,-64.5,87,-63.5</points>
<connection>
<GID>17</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>92.5,-64.5,92.5,-63.5</points>
<connection>
<GID>19</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>98,-64.5,98,-63.5</points>
<connection>
<GID>21</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>103.5,-64.5,103.5,-63.5</points>
<connection>
<GID>23</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>109,-66,109,-63.5</points>
<connection>
<GID>25</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>114.5,-64.5,114.5,-63.5</points>
<connection>
<GID>27</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>120,-64.5,120,-63.5</points>
<connection>
<GID>28</GID>
<name>SEL_0</name></connection>
<intersection>-63.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-14.5,3,-14</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-14,3,-14</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,2.5,-3,4</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,2.5,-1,4</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,0.5,1.5,2</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,0.5,3.5,2</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>5.5,-2,5.5,2</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-62.5,77.5,-62.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-62.5,79.5,-62.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-14.5,7,-9.5</points>
<connection>
<GID>8</GID>
<name>IN_4</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-14.5,8,-14.5</points>
<connection>
<GID>8</GID>
<name>IN_5</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-14.5,9,-9.5</points>
<connection>
<GID>8</GID>
<name>IN_6</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-14.5,11.5,-14.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-9,12,-3.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17.5,-14.5,17.5,-9</points>
<intersection>-14.5 3</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12,-9,17.5,-9</points>
<intersection>12 0</intersection>
<intersection>17.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-14.5,18,-14.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>17.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-8,16.5,-5.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>19,-14.5,19,-8</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-8,19,-8</points>
<intersection>16.5 0</intersection>
<intersection>19 1</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-14.5,20,-5</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-14.5,17,-14</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14,-14,17,-14</points>
<intersection>14 3</intersection>
<intersection>17 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-14,14,-13.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,2.5,11,3.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,2.5,13,4.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,0.5,15.5,3.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,0.5,17.5,1.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-1,20,2.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>2.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,2.5,20.5,2.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-14.5,21,-9.5</points>
<connection>
<GID>59</GID>
<name>IN_4</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-14.5,22,-14.5</points>
<connection>
<GID>59</GID>
<name>IN_5</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-14.5,23,-9.5</points>
<connection>
<GID>59</GID>
<name>IN_6</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-14.5,24,-14.5</points>
<connection>
<GID>59</GID>
<name>IN_7</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-9.5,25.5,-4</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,-15,31,-9.5</points>
<intersection>-15 3</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-9.5,31,-9.5</points>
<intersection>25.5 0</intersection>
<intersection>31 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-15,31.5,-15</points>
<intersection>31 1</intersection>
<intersection>31.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31.5,-15.5,31.5,-15</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-15 3</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-8.5,30,-6</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32.5,-15.5,32.5,-8.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,-8.5,32.5,-8.5</points>
<intersection>30 0</intersection>
<intersection>32.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-15.5,33.5,-5.5</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-15.5,30.5,-14.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-14.5,30.5,-14.5</points>
<intersection>27.5 4</intersection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-14.5,27.5,-14</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>24.5,2,24.5,4.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>26.5,2,26.5,4</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>29,-1.19249e-008,29,2</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>31,1.19249e-008,31,1</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>33.5,-1.5,33.5,-1</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-15.5,34.5,-10</points>
<connection>
<GID>73</GID>
<name>IN_4</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-15.5,35.5,-15</points>
<connection>
<GID>73</GID>
<name>IN_5</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-15.5,36.5,-10</points>
<connection>
<GID>73</GID>
<name>IN_6</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-15.5,37.5,-15</points>
<connection>
<GID>73</GID>
<name>IN_7</name></connection>
<connection>
<GID>86</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-9.5,39.5,-4</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>-9.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45,-15,45,-9.5</points>
<intersection>-15 3</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-9.5,45,-9.5</points>
<intersection>39.5 0</intersection>
<intersection>45 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45,-15,45.5,-15</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>45 1</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-8.5,44,-6</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46.5,-15,46.5,-8.5</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44,-8.5,46.5,-8.5</points>
<intersection>44 0</intersection>
<intersection>46.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-15,47.5,-5</points>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-15,44.5,-14.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-14.5,44.5,-14.5</points>
<intersection>41.5 6</intersection>
<intersection>44.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>41.5,-14.5,41.5,-14</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,2,38.5,3.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,2,40.5,3</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-1.19249e-008,43,0.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,1.19249e-008,45,1</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-1,47.5,-0.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-15,48.5,-10.5</points>
<connection>
<GID>87</GID>
<name>IN_4</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-15,50,-15</points>
<connection>
<GID>87</GID>
<name>IN_5</name></connection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-15,50,-12.5</points>
<intersection>-15 1</intersection>
<intersection>-12.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50,-12.5,50.5,-12.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>50 4</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-14,52,-6.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-14,52,-14</points>
<intersection>50.5 3</intersection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-15,50.5,-14</points>
<connection>
<GID>87</GID>
<name>IN_6</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-15,53.5,-13.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-15,53.5,-15</points>
<connection>
<GID>87</GID>
<name>IN_7</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-14.5,56,-7</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-14.5,57.5,-14.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-62.5,83.5,-62.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-62.5,85.5,-62.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-62.5,89,-62</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-62.5,91,-62</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-62.5,94.5,-62.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-62.5,97,-62.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-62.5,100,-62.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-62.5,102,-62.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-64,105.5,-62.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-64,107.5,-62.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-62.5,111,-62.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-62.5,113,-62.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-62.5,116.5,-62.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-14.5,58,-11.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-14.5,58.5,-14.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-14.5,59.5,-7</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<connection>
<GID>119</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-14.5,60.5,-13</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<connection>
<GID>120</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-14.5,61.5,-9</points>
<connection>
<GID>10</GID>
<name>IN_4</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-62.5,119,-62.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-14.5,63.5,-10</points>
<connection>
<GID>10</GID>
<name>IN_6</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-14.5,64.5,-14</points>
<connection>
<GID>10</GID>
<name>IN_7</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-14,69.5,-6.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-14,71,-14</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-14,71.5,-11</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-14,72,-14</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-14,72.5,-6.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-14 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,-14,73,-14</points>
<connection>
<GID>125</GID>
<name>IN_2</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-14,74,-12.5</points>
<connection>
<GID>125</GID>
<name>IN_3</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-14,75,-8.5</points>
<connection>
<GID>125</GID>
<name>IN_4</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,87,80,89</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-14,77,-9.5</points>
<connection>
<GID>125</GID>
<name>IN_6</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-14,78,-13.5</points>
<connection>
<GID>125</GID>
<name>IN_7</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-13.5,82,-6</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-13.5,83.5,-13.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-13.5,84,-10.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-13.5,84.5,-13.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-13.5,85.5,-6</points>
<connection>
<GID>134</GID>
<name>IN_2</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-13.5,86.5,-12</points>
<connection>
<GID>134</GID>
<name>IN_3</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-13.5,87.5,-8</points>
<connection>
<GID>134</GID>
<name>IN_4</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,87,82,89</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,57,-19,59</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-13.5,93,-11.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-13.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>90.5,-13.5,93,-13.5</points>
<connection>
<GID>134</GID>
<name>IN_7</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-13.5,96,-6</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-13.5,97.5,-13.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-13.5,98,-10.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-13.5,98.5,-13.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-13.5,99.5,-6</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-13.5,100.5,-12</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-13.5,101.5,-8</points>
<connection>
<GID>143</GID>
<name>IN_4</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,57,-17,59</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-13.5,103.5,-9</points>
<connection>
<GID>143</GID>
<name>IN_6</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-13.5,106.5,-10</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-13.5,106.5,-13.5</points>
<connection>
<GID>143</GID>
<name>IN_7</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,57,-14.5,59</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,57,-12.5,59</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,57,-10,59</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,57,-8,59</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,57,-5,59</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,57,-3,59</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35,-109.5,-31,-109.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>153</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-35.5,-118.5,-30.5,-118.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-30.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-30.5,-120,-30.5,-118.5</points>
<connection>
<GID>155</GID>
<name>clock</name></connection>
<intersection>-118.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,5,76,6</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,5.5,89,6.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,4.5,102.5,6</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,4,62.5,5.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-14.5,62.5,0</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-14,76,1</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-6,89,1.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>88.5,-13.5,88.5,-6</points>
<connection>
<GID>134</GID>
<name>IN_5</name></connection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-6,89,-6</points>
<intersection>88.5 1</intersection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-13.5,102.5,0.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-13.5,89.5,-11</points>
<connection>
<GID>134</GID>
<name>IN_6</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>90,-11,90,-9</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-11,90,-11</points>
<intersection>89.5 0</intersection>
<intersection>90 1</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-35,6.5,-20.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>-35 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48,-38,48,-35</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-35,48,-35</points>
<intersection>6.5 0</intersection>
<intersection>48 1</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-131,-31,-130.5</points>
<connection>
<GID>157</GID>
<name>clock</name></connection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-130.5,-31,-130.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-28,48,-21</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-38,53,-28</points>
<intersection>-38 3</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48,-28,53,-28</points>
<intersection>48 0</intersection>
<intersection>53 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51,-38,53,-38</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>53 1</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-30,34,-21.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-38,50,-30</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34,-30,50,-30</points>
<intersection>34 0</intersection>
<intersection>50 1</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-38,49,-31.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-31.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,-31.5,20.5,-20.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-31.5,49,-31.5</points>
<intersection>20.5 1</intersection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-30,101,-19.5</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58,-38,58,-30</points>
<connection>
<GID>20</GID>
<name>IN_B_0</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,-30,101,-30</points>
<intersection>58 1</intersection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-28.5,87,-19.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57,-38,57,-28.5</points>
<connection>
<GID>20</GID>
<name>IN_B_1</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-28.5,87,-28.5</points>
<intersection>57 1</intersection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-38,56,-33</points>
<connection>
<GID>20</GID>
<name>IN_B_2</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>74.5,-33,74.5,-20</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56,-33,74.5,-33</points>
<intersection>56 0</intersection>
<intersection>74.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-38,55.5,-22.5</points>
<intersection>-38 5</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>55.5,-22.5,61,-22.5</points>
<intersection>55.5 0</intersection>
<intersection>61 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>61,-22.5,61,-20.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>55,-38,55.5,-38</points>
<connection>
<GID>20</GID>
<name>IN_B_3</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-44,120,-23</points>
<intersection>-44 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-23,120,-23</points>
<intersection>-2.5 22</intersection>
<intersection>15.5 4</intersection>
<intersection>29 7</intersection>
<intersection>43.5 10</intersection>
<intersection>55 12</intersection>
<intersection>69.5 14</intersection>
<intersection>82.5 16</intersection>
<intersection>96 20</intersection>
<intersection>117.5 18</intersection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-44,120,-44</points>
<intersection>93.5 3</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>93.5,-44,93.5,-40.5</points>
<connection>
<GID>18</GID>
<name>SEL_2</name></connection>
<intersection>-44 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>15.5,-23,15.5,-16.5</points>
<intersection>-23 1</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>12,-16.5,15.5,-16.5</points>
<connection>
<GID>8</GID>
<name>SEL_2</name></connection>
<intersection>15.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-23,29,-16.5</points>
<intersection>-23 1</intersection>
<intersection>-16.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>26,-16.5,29,-16.5</points>
<connection>
<GID>59</GID>
<name>SEL_2</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>43.5,-23,43.5,-17.5</points>
<intersection>-23 1</intersection>
<intersection>-17.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>39.5,-17.5,43.5,-17.5</points>
<connection>
<GID>73</GID>
<name>SEL_2</name></connection>
<intersection>43.5 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>55,-23,55,-17</points>
<intersection>-23 1</intersection>
<intersection>-17 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>53.5,-17,55,-17</points>
<connection>
<GID>87</GID>
<name>SEL_2</name></connection>
<intersection>55 12</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>69.5,-23,69.5,-16.5</points>
<intersection>-23 1</intersection>
<intersection>-16.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>66.5,-16.5,69.5,-16.5</points>
<connection>
<GID>10</GID>
<name>SEL_2</name></connection>
<intersection>69.5 14</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>82.5,-23,82.5,-16</points>
<intersection>-23 1</intersection>
<intersection>-16 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>80,-16,82.5,-16</points>
<connection>
<GID>125</GID>
<name>SEL_2</name></connection>
<intersection>82.5 16</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>117.5,-23,117.5,-15.5</points>
<intersection>-23 1</intersection>
<intersection>-15.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>106.5,-15.5,117.5,-15.5</points>
<connection>
<GID>143</GID>
<name>SEL_2</name></connection>
<intersection>117.5 18</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>96,-23,96,-15.5</points>
<intersection>-23 1</intersection>
<intersection>-15.5 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>92.5,-15.5,96,-15.5</points>
<connection>
<GID>134</GID>
<name>SEL_2</name></connection>
<intersection>96 20</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-2.5,-24.5,-2.5,-23</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-110,-6,-109</points>
<intersection>-110 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-110,-6,-110</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-109,-5.5,-109</points>
<connection>
<GID>161</GID>
<name>clock</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-46,116,-26</points>
<intersection>-46 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-26,116,-26</points>
<intersection>-2.5 10</intersection>
<intersection>14.5 4</intersection>
<intersection>27.5 7</intersection>
<intersection>42.5 11</intersection>
<intersection>54.5 13</intersection>
<intersection>68 16</intersection>
<intersection>82 18</intersection>
<intersection>95 23</intersection>
<intersection>114.5 21</intersection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-46,116,-46</points>
<intersection>92.5 3</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-46,92.5,-40.5</points>
<connection>
<GID>18</GID>
<name>SEL_1</name></connection>
<intersection>-46 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>14.5,-26,14.5,-17.5</points>
<intersection>-26 1</intersection>
<intersection>-17.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>12,-17.5,14.5,-17.5</points>
<connection>
<GID>8</GID>
<name>SEL_1</name></connection>
<intersection>14.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>27.5,-26,27.5,-17.5</points>
<intersection>-26 1</intersection>
<intersection>-17.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>26,-17.5,27.5,-17.5</points>
<connection>
<GID>59</GID>
<name>SEL_1</name></connection>
<intersection>27.5 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-2.5,-26.5,-2.5,-26</points>
<intersection>-26.5 15</intersection>
<intersection>-26 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>42.5,-26,42.5,-18.5</points>
<intersection>-26 1</intersection>
<intersection>-18.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>39.5,-18.5,42.5,-18.5</points>
<connection>
<GID>73</GID>
<name>SEL_1</name></connection>
<intersection>42.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>54.5,-26,54.5,-18</points>
<intersection>-26 1</intersection>
<intersection>-18 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>53.5,-18,54.5,-18</points>
<connection>
<GID>87</GID>
<name>SEL_1</name></connection>
<intersection>54.5 13</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-8,-26.5,-2.5,-26.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-2.5 10</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>68,-26,68,-17.5</points>
<intersection>-26 1</intersection>
<intersection>-17.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>66.5,-17.5,68,-17.5</points>
<connection>
<GID>10</GID>
<name>SEL_1</name></connection>
<intersection>68 16</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>82,-26,82,-17</points>
<intersection>-26 1</intersection>
<intersection>-17 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>80,-17,82,-17</points>
<connection>
<GID>125</GID>
<name>SEL_1</name></connection>
<intersection>82 18</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>114.5,-26,114.5,-16.5</points>
<intersection>-26 1</intersection>
<intersection>-16.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>106.5,-16.5,114.5,-16.5</points>
<connection>
<GID>143</GID>
<name>SEL_1</name></connection>
<intersection>114.5 21</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>95,-26,95,-16.5</points>
<intersection>-26 1</intersection>
<intersection>-16.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>92.5,-16.5,95,-16.5</points>
<connection>
<GID>134</GID>
<name>SEL_1</name></connection>
<intersection>95 23</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-48.5,114,-27</points>
<intersection>-48.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-27,114,-27</points>
<intersection>-2.5 6</intersection>
<intersection>13.5 4</intersection>
<intersection>26 11</intersection>
<intersection>41 7</intersection>
<intersection>53.5 9</intersection>
<intersection>66.5 10</intersection>
<intersection>80 12</intersection>
<intersection>93 15</intersection>
<intersection>112 13</intersection>
<intersection>114 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-48.5,114,-48.5</points>
<intersection>91.5 3</intersection>
<intersection>114 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-48.5,91.5,-40.5</points>
<connection>
<GID>18</GID>
<name>SEL_0</name></connection>
<intersection>-48.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>13.5,-27,13.5,-18.5</points>
<intersection>-27 1</intersection>
<intersection>-18.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>12,-18.5,13.5,-18.5</points>
<connection>
<GID>8</GID>
<name>SEL_0</name></connection>
<intersection>13.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-2.5,-31,-2.5,-27</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>41,-27,41,-19.5</points>
<intersection>-27 1</intersection>
<intersection>-19.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>39.5,-19.5,41,-19.5</points>
<connection>
<GID>73</GID>
<name>SEL_0</name></connection>
<intersection>41 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>53.5,-27,53.5,-19</points>
<connection>
<GID>87</GID>
<name>SEL_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>66.5,-27,66.5,-18.5</points>
<connection>
<GID>10</GID>
<name>SEL_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>26,-27,26,-18.5</points>
<connection>
<GID>59</GID>
<name>SEL_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>80,-27,80,-18</points>
<connection>
<GID>125</GID>
<name>SEL_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>112,-27,112,-17.5</points>
<intersection>-27 1</intersection>
<intersection>-17.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>106.5,-17.5,112,-17.5</points>
<connection>
<GID>143</GID>
<name>SEL_0</name></connection>
<intersection>112 13</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>93,-27,93,-17.5</points>
<intersection>-27 1</intersection>
<intersection>-17.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>92.5,-17.5,93,-17.5</points>
<connection>
<GID>134</GID>
<name>SEL_0</name></connection>
<intersection>93 15</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-41,75,-35</points>
<intersection>-41 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-41,75,-41</points>
<connection>
<GID>20</GID>
<name>carry_in</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-35,89.5,-35</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-47.5,-10.5,-44</points>
<intersection>-47.5 5</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,-44,-7.5,-44</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-47.5,-10.5,-47.5</points>
<connection>
<GID>175</GID>
<name>OUT_3</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-49,-8.5,-49</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-10.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-10.5,-49.5,-10.5,-49</points>
<intersection>-49.5 6</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-12.5,-49.5,-10.5,-49.5</points>
<connection>
<GID>175</GID>
<name>OUT_2</name></connection>
<intersection>-10.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12.5,-51.5,-6.5,-51.5</points>
<connection>
<GID>175</GID>
<name>OUT_1</name></connection>
<intersection>-6.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-6.5,-52,-6.5,-51.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-55.5,-10.5,-53.5</points>
<intersection>-55.5 1</intersection>
<intersection>-53.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,-55.5,-9,-55.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-53.5,-10.5,-53.5</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-47,12,-44</points>
<intersection>-47 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-44,15,-44</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-47,12,-47</points>
<connection>
<GID>191</GID>
<name>OUT_3</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-49,14,-49</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<connection>
<GID>191</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-51.5,12,-51</points>
<intersection>-51.5 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-51.5,16,-51.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-51,12,-51</points>
<connection>
<GID>191</GID>
<name>OUT_1</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-55.5,12,-53</points>
<intersection>-55.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-55.5,13.5,-55.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-53,12,-53</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-47,32.5,-44</points>
<intersection>-47 6</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-44,35.5,-44</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>30,-47,32.5,-47</points>
<connection>
<GID>196</GID>
<name>OUT_3</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>30,-49,34.5,-49</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>196</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-51,36.5,-51</points>
<connection>
<GID>196</GID>
<name>OUT_1</name></connection>
<intersection>36.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>36.5,-51.5,36.5,-51</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-55.5,32.5,-53</points>
<intersection>-55.5 1</intersection>
<intersection>-53 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-55.5,34,-55.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>30,-53,32.5,-53</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-69.5,26,-67</points>
<intersection>-69.5 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-67,26,-67</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-69.5,28.5,-69.5</points>
<connection>
<GID>185</GID>
<name>IN_3</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-70.5,28.5,-70.5</points>
<connection>
<GID>185</GID>
<name>IN_2</name></connection>
<intersection>21.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>21.5,-70.5,21.5,-70</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-71.5,28.5,-71.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<connection>
<GID>204</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-74.5,27,-74.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>27 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>27,-74.5,27,-72.5</points>
<intersection>-74.5 1</intersection>
<intersection>-72.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>27,-72.5,28.5,-72.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>27 5</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-68.5,52.5,-66</points>
<intersection>-68.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-66,52.5,-66</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-68.5,55,-68.5</points>
<connection>
<GID>210</GID>
<name>IN_3</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-69.5,55,-69.5</points>
<connection>
<GID>210</GID>
<name>IN_2</name></connection>
<intersection>48 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>48,-69.5,48,-69</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>-69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-70.5,55,-70.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-73.5,53.5,-73.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>53.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53.5,-73.5,53.5,-71.5</points>
<intersection>-73.5 1</intersection>
<intersection>-71.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>53.5,-71.5,55,-71.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>53.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-49.5,53,-46</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-46,53.5,-46</points>
<connection>
<GID>20</GID>
<name>OUT_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-50.5,55.5,-46</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-46,55.5,-46</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-52,50.5,-47.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-47.5,52.5,-47.5</points>
<intersection>50.5 0</intersection>
<intersection>52.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>52.5,-47.5,52.5,-46</points>
<connection>
<GID>20</GID>
<name>OUT_2</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-50.5,46.5,-49</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-49,51.5,-49</points>
<intersection>46.5 0</intersection>
<intersection>51.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>51.5,-49,51.5,-46</points>
<connection>
<GID>20</GID>
<name>OUT_3</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-7,-120.5,-5.5,-120.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-5.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-5.5,-120.5,-5.5,-120</points>
<connection>
<GID>167</GID>
<name>clock</name></connection>
<intersection>-120.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-131.5,-6,-131</points>
<connection>
<GID>170</GID>
<name>clock</name></connection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-131.5,-6,-131.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-108.5,20.5,-108.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>20,-119,21,-119</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<connection>
<GID>180</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-130.5,20.5,-130</points>
<connection>
<GID>183</GID>
<name>clock</name></connection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-130.5,20.5,-130.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-108,49.5,-107.5</points>
<connection>
<GID>211</GID>
<name>clock</name></connection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-108,49.5,-108</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>47,-118,50,-118</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-129,49.5,-128.5</points>
<connection>
<GID>219</GID>
<name>clock</name></connection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-128.5,49.5,-128.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-107,81,-106.5</points>
<connection>
<GID>254</GID>
<name>clock</name></connection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-107,81,-107</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>78.5,-117,81.5,-117</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<connection>
<GID>261</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-128,81,-128</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<connection>
<GID>265</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-106,108,-106</points>
<connection>
<GID>273</GID>
<name>clock</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>108,-116.5,108.5,-116.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<connection>
<GID>277</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-127.5,108,-127.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-105.5,134.5,-105</points>
<connection>
<GID>286</GID>
<name>clock</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,-105,134.5,-105</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-116,133.5,-115</points>
<intersection>-116 9</intersection>
<intersection>-115 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>133.5,-116,135,-116</points>
<connection>
<GID>288</GID>
<name>clock</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>132.5,-115,133.5,-115</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-127,134.5,-126.5</points>
<connection>
<GID>290</GID>
<name>clock</name></connection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-126.5,134.5,-126.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160.5,-106.5,162.5,-106.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<connection>
<GID>294</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>161,-117,162.5,-117</points>
<connection>
<GID>296</GID>
<name>clock</name></connection>
<intersection>161 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>161,-117,161,-115.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-117 5</intersection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-128,161,-126.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-128,163,-128</points>
<connection>
<GID>298</GID>
<name>clock</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159,-153,161.5,-153</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>161.5,-163.5,162,-163.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<connection>
<GID>304</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,44,1,47.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>0.5,47.5,0.5,51</points>
<intersection>47.5 2</intersection>
<intersection>51 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0.5,47.5,1,47.5</points>
<intersection>0.5 1</intersection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4,51,0.5,51</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>0.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,44,0,47.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-9,47.5,-9,51</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-9,47.5,0,47.5</points>
<intersection>-9 1</intersection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,46.5,-13.5,51</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1,44,-1,46.5</points>
<connection>
<GID>106</GID>
<name>IN_2</name></connection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,46.5,-1,46.5</points>
<intersection>-13.5 0</intersection>
<intersection>-1 1</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,45,-18,51</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-2,44,-2,45</points>
<connection>
<GID>106</GID>
<name>IN_3</name></connection>
<intersection>45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-18,45,-2,45</points>
<intersection>-18 0</intersection>
<intersection>-2 1</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,77,6,79</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<connection>
<GID>221</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,77,8,79</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,77,10.5,79</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,77,12.5,79</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,77,15,79</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,77,17,79</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,77,20,79</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,77,22,79</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,64,26,67.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>67.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,67.5,25.5,71</points>
<intersection>67.5 2</intersection>
<intersection>71 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25.5,67.5,26,67.5</points>
<intersection>25.5 1</intersection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21,71,25.5,71</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<intersection>25.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,64,25,67.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>67.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>16,67.5,16,71</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<intersection>67.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16,67.5,25,67.5</points>
<intersection>16 1</intersection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,66.5,11.5,71</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>24,64,24,66.5</points>
<connection>
<GID>228</GID>
<name>IN_2</name></connection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,66.5,24,66.5</points>
<intersection>11.5 0</intersection>
<intersection>24 1</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,65,7,71</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>65 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>23,64,23,65</points>
<connection>
<GID>228</GID>
<name>IN_3</name></connection>
<intersection>65 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,65,23,65</points>
<intersection>7 0</intersection>
<intersection>23 1</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,88.5,34,90.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,88.5,36,90.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,88.5,38.5,90.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,88.5,40.5,90.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>238</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,88.5,43,90.5</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,88.5,45,90.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,88.5,48,90.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,88.5,50,90.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,75.5,54,79</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53.5,79,53.5,82.5</points>
<intersection>79 2</intersection>
<intersection>82.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53.5,79,54,79</points>
<intersection>53.5 1</intersection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>49,82.5,53.5,82.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>53.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,75.5,53,79</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,79,44,82.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44,79,53,79</points>
<intersection>44 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,78,39.5,82.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,75.5,52,78</points>
<connection>
<GID>241</GID>
<name>IN_2</name></connection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,78,52,78</points>
<intersection>39.5 0</intersection>
<intersection>52 1</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,76.5,35,82.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>76.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51,75.5,51,76.5</points>
<connection>
<GID>241</GID>
<name>IN_3</name></connection>
<intersection>76.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,76.5,51,76.5</points>
<intersection>35 0</intersection>
<intersection>51 1</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-174.5,161.5,-174</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<intersection>-174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,-174,161.5,-174</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-153,134,-153</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>310</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,92.5,62,94.5</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,92.5,64,94.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<connection>
<GID>251</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,92.5,66.5,94.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<connection>
<GID>253</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,92.5,68.5,94.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,92.5,71.5,94.5</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,92.5,73.5,94.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>132,-163.5,134.5,-163.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<connection>
<GID>312</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132,-174.5,134,-174.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>314</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-154,108,-152.5</points>
<connection>
<GID>318</GID>
<name>clock</name></connection>
<intersection>-154 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-154,108,-154</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>106.5,-163,108.5,-163</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<connection>
<GID>320</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,77.5,72.5,86.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>77.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>61,75.5,61,77.5</points>
<connection>
<GID>241</GID>
<name>IN_B_0</name></connection>
<intersection>77.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,77.5,72.5,77.5</points>
<intersection>61 1</intersection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,81,63,86.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59,75.5,59,81</points>
<connection>
<GID>241</GID>
<name>IN_B_2</name></connection>
<intersection>81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,81,63,81</points>
<intersection>59 1</intersection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,79.5,67.5,86.5</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<intersection>79.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60,75.5,60,79.5</points>
<connection>
<GID>241</GID>
<name>IN_B_1</name></connection>
<intersection>79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,79.5,67.5,79.5</points>
<intersection>60 1</intersection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-174,108,-174</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>322</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,44,5,61</points>
<connection>
<GID>106</GID>
<name>IN_B_3</name></connection>
<intersection>61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,61,20,61</points>
<connection>
<GID>228</GID>
<name>carry_out</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,44,6,56</points>
<connection>
<GID>106</GID>
<name>IN_B_2</name></connection>
<intersection>56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>6,56,26.5,56</points>
<connection>
<GID>228</GID>
<name>OUT_3</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,54,27.5,56</points>
<connection>
<GID>228</GID>
<name>OUT_2</name></connection>
<intersection>54 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>7,44,7,54</points>
<connection>
<GID>106</GID>
<name>IN_B_1</name></connection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,54,27.5,54</points>
<intersection>7 1</intersection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,50,28.5,56</points>
<connection>
<GID>228</GID>
<name>OUT_1</name></connection>
<intersection>50 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8,44,8,50</points>
<connection>
<GID>106</GID>
<name>IN_B_0</name></connection>
<intersection>50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,50,28.5,50</points>
<intersection>8 1</intersection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,41,12,41</points>
<connection>
<GID>106</GID>
<name>carry_in</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,30,6,36</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,36,6,36</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,30,3.5,36</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,25,2,36</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,36,2.5,36</points>
<connection>
<GID>106</GID>
<name>OUT_2</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,27,-1,36</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,36,1.5,36</points>
<connection>
<GID>106</GID>
<name>OUT_3</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,41,-5,41</points>
<connection>
<GID>106</GID>
<name>carry_out</name></connection>
<intersection>-6 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-6,28,-6,41</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,50.5,30,56</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,56,30,56</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,64,30,72.5</points>
<connection>
<GID>228</GID>
<name>IN_B_3</name></connection>
<intersection>72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,72.5,48,72.5</points>
<connection>
<GID>241</GID>
<name>carry_out</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,66.5,54.5,67.5</points>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<intersection>66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,64,31,66.5</points>
<connection>
<GID>228</GID>
<name>IN_B_2</name></connection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31,66.5,54.5,66.5</points>
<intersection>31 1</intersection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,65.5,55.5,67.5</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<intersection>65.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32,64,32,65.5</points>
<connection>
<GID>228</GID>
<name>IN_B_1</name></connection>
<intersection>65.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,65.5,55.5,65.5</points>
<intersection>32 1</intersection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,64.5,56.5,67.5</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<intersection>64.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33,64,33,64.5</points>
<connection>
<GID>228</GID>
<name>IN_B_0</name></connection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,64.5,56.5,64.5</points>
<intersection>33 1</intersection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,65.5,57.5,67.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<connection>
<GID>274</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,72.5,64,72.5</points>
<connection>
<GID>241</GID>
<name>carry_in</name></connection>
<connection>
<GID>276</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,80.5,81,81</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,75.5,58,82.5</points>
<connection>
<GID>241</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,60.5,36,61</points>
<connection>
<GID>228</GID>
<name>carry_in</name></connection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,60.5,38,60.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-153,80,-153</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>73.5,-164.5,80.5,-164.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>80.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>80.5,-164.5,80.5,-163.5</points>
<connection>
<GID>328</GID>
<name>clock</name></connection>
<intersection>-164.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-174.5,79.5,-174.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<connection>
<GID>330</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-155,21,-154</points>
<connection>
<GID>334</GID>
<name>clock</name></connection>
<intersection>-154 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-154,21,-154</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>18.5,-164,21.5,-164</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>21.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>21.5,-165,21.5,-164</points>
<connection>
<GID>336</GID>
<name>clock</name></connection>
<intersection>-164 5</intersection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-176,21,-176</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-153.5,49.5,-153.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>47,-164,50,-164</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>344</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-175.5,49.5,-175</points>
<connection>
<GID>346</GID>
<name>clock</name></connection>
<intersection>-175.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-175.5,49.5,-175.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-154,-6,-154</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>350</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-7.5,-164.5,-5.5,-164.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>352</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-175.5,-6,-175</points>
<connection>
<GID>354</GID>
<name>clock</name></connection>
<intersection>-175 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-175,-6,-175</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-154.5,-31,-154</points>
<connection>
<GID>358</GID>
<name>clock</name></connection>
<intersection>-154.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-154.5,-31,-154.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-32.5,-164.5,-30.5,-164.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<connection>
<GID>360</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34,-175.5,-31,-175.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<connection>
<GID>362</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-129,-62,-100.5</points>
<connection>
<GID>366</GID>
<name>OUT_7</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-62,-100.5,165.5,-100.5</points>
<connection>
<GID>286</GID>
<name>set</name></connection>
<intersection>-62 0</intersection>
<intersection>-28 13</intersection>
<intersection>-2.5 12</intersection>
<intersection>23.5 5</intersection>
<intersection>52.5 14</intersection>
<intersection>84 20</intersection>
<intersection>111 15</intersection>
<intersection>165.5 19</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23.5,-103.5,23.5,-100.5</points>
<connection>
<GID>178</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-2.5,-104,-2.5,-100.5</points>
<connection>
<GID>161</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-28,-104.5,-28,-100.5</points>
<connection>
<GID>153</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>52.5,-102.5,52.5,-100.5</points>
<connection>
<GID>211</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-101,111,-100.5</points>
<connection>
<GID>273</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>165.5,-101.5,165.5,-100.5</points>
<connection>
<GID>294</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>84,-101.5,84,-100.5</points>
<connection>
<GID>254</GID>
<name>set</name></connection>
<intersection>-100.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-138,161.5,-137.5</points>
<intersection>-138 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-138,162.5,-138</points>
<connection>
<GID>300</GID>
<name>clock</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160.5,-137.5,161.5,-137.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-185.5,160,-185</points>
<intersection>-185.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-185,161.5,-185</points>
<connection>
<GID>308</GID>
<name>clock</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>159,-185.5,160,-185.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-185,132,-184</points>
<intersection>-185 1</intersection>
<intersection>-184 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-185,134,-185</points>
<connection>
<GID>316</GID>
<name>clock</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130.5,-184,132,-184</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,-141.5,-31,-141.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-186,-32.5,-184.5</points>
<intersection>-186 1</intersection>
<intersection>-184.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-186,-31,-186</points>
<connection>
<GID>364</GID>
<name>clock</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-184.5,-32.5,-184.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-186,-9.5,-185.5</points>
<intersection>-186 1</intersection>
<intersection>-185.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-186,-6,-186</points>
<connection>
<GID>356</GID>
<name>clock</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-185.5,-9.5,-185.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-186.5,21,-186.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-185.5,48.5,-185</points>
<intersection>-185.5 1</intersection>
<intersection>-185 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-185.5,49.5,-185.5</points>
<connection>
<GID>348</GID>
<name>clock</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-185,48.5,-185</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-185.5,78.5,-185</points>
<intersection>-185.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-185,79.5,-185</points>
<connection>
<GID>332</GID>
<name>clock</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-185.5,78.5,-185.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-185,106.5,-184.5</points>
<intersection>-185 2</intersection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-184.5,108,-184.5</points>
<connection>
<GID>324</GID>
<name>clock</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-185,106.5,-185</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-142,-7.5,-141.5</points>
<intersection>-142 2</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-141.5,-6,-141.5</points>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-9,-142,-7.5,-142</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-140.5,20.5,-140.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>186</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-140,47.5,-139.5</points>
<intersection>-140 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-139.5,49,-139.5</points>
<connection>
<GID>247</GID>
<name>clock</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-140,47.5,-140</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-139,81,-139</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>81 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-139,81,-138.5</points>
<connection>
<GID>269</GID>
<name>clock</name></connection>
<intersection>-139 1</intersection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-138.5,106,-138</points>
<intersection>-138.5 2</intersection>
<intersection>-138 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-138,108,-138</points>
<connection>
<GID>284</GID>
<name>clock</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-138.5,106,-138.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-137.5,133,-137</points>
<intersection>-137.5 1</intersection>
<intersection>-137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-137.5,134.5,-137.5</points>
<connection>
<GID>292</GID>
<name>clock</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-137,133,-137</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-130,-61.5,-115</points>
<intersection>-130 1</intersection>
<intersection>-115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-130,-61.5,-130</points>
<connection>
<GID>366</GID>
<name>OUT_6</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-61.5,-115,24,-115</points>
<connection>
<GID>167</GID>
<name>set</name></connection>
<connection>
<GID>155</GID>
<name>set</name></connection>
<intersection>-61.5 0</intersection>
<intersection>24 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,-115,24,-113</points>
<connection>
<GID>180</GID>
<name>set</name></connection>
<intersection>-115 2</intersection>
<intersection>-113 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>24,-113,84.5,-113</points>
<connection>
<GID>217</GID>
<name>set</name></connection>
<intersection>24 4</intersection>
<intersection>84.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>84.5,-113,84.5,-111.5</points>
<connection>
<GID>261</GID>
<name>set</name></connection>
<intersection>-113 5</intersection>
<intersection>-111.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-111.5,165.5,-111.5</points>
<connection>
<GID>277</GID>
<name>set</name></connection>
<intersection>84.5 6</intersection>
<intersection>138 13</intersection>
<intersection>165.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>165.5,-112,165.5,-111.5</points>
<connection>
<GID>296</GID>
<name>set</name></connection>
<intersection>-111.5 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>138,-111.5,138,-111</points>
<connection>
<GID>288</GID>
<name>set</name></connection>
<intersection>-111.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61,-130.5,-61,-126</points>
<intersection>-130.5 1</intersection>
<intersection>-126 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-130.5,-61,-130.5</points>
<intersection>-62 2</intersection>
<intersection>-61 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-62,-131,-62,-130.5</points>
<connection>
<GID>366</GID>
<name>OUT_5</name></connection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-61,-126,23.5,-126</points>
<connection>
<GID>170</GID>
<name>set</name></connection>
<connection>
<GID>157</GID>
<name>set</name></connection>
<intersection>-61 0</intersection>
<intersection>23.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23.5,-126,23.5,-124</points>
<connection>
<GID>183</GID>
<name>set</name></connection>
<intersection>-126 3</intersection>
<intersection>-124 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>23.5,-124,84,-124</points>
<connection>
<GID>219</GID>
<name>set</name></connection>
<intersection>23.5 5</intersection>
<intersection>84 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>84,-124,84,-122.5</points>
<connection>
<GID>265</GID>
<name>set</name></connection>
<intersection>-124 6</intersection>
<intersection>-122.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>84,-122.5,166,-122.5</points>
<connection>
<GID>281</GID>
<name>set</name></connection>
<intersection>84 7</intersection>
<intersection>137.5 9</intersection>
<intersection>166 10</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>137.5,-122.5,137.5,-122</points>
<connection>
<GID>290</GID>
<name>set</name></connection>
<intersection>-122.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>166,-123,166,-122.5</points>
<connection>
<GID>298</GID>
<name>set</name></connection>
<intersection>-122.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-136.5,-58,-132</points>
<intersection>-136.5 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-132,-58,-132</points>
<connection>
<GID>366</GID>
<name>OUT_4</name></connection>
<intersection>-58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-58,-136.5,23.5,-136.5</points>
<connection>
<GID>176</GID>
<name>set</name></connection>
<connection>
<GID>159</GID>
<name>set</name></connection>
<intersection>-58 0</intersection>
<intersection>23.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-136.5,23.5,-134.5</points>
<connection>
<GID>186</GID>
<name>set</name></connection>
<intersection>-136.5 2</intersection>
<intersection>-134.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23.5,-134.5,84,-134.5</points>
<connection>
<GID>247</GID>
<name>set</name></connection>
<intersection>23.5 4</intersection>
<intersection>84 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>84,-134.5,84,-133</points>
<connection>
<GID>269</GID>
<name>set</name></connection>
<intersection>-134.5 5</intersection>
<intersection>-133 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>84,-133,165.5,-133</points>
<connection>
<GID>300</GID>
<name>set</name></connection>
<connection>
<GID>284</GID>
<name>set</name></connection>
<intersection>84 6</intersection>
<intersection>137.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>137.5,-133,137.5,-132.5</points>
<connection>
<GID>292</GID>
<name>set</name></connection>
<intersection>-133 7</intersection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-148.5,-57,-133</points>
<intersection>-148.5 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-133,-57,-133</points>
<connection>
<GID>366</GID>
<name>OUT_3</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-148.5,52.5,-148.5</points>
<intersection>-57 0</intersection>
<intersection>-28 8</intersection>
<intersection>-3 9</intersection>
<intersection>24 4</intersection>
<intersection>52.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,-150,24,-148.5</points>
<connection>
<GID>334</GID>
<name>set</name></connection>
<intersection>-148.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>52.5,-148.5,52.5,-148</points>
<connection>
<GID>342</GID>
<name>set</name></connection>
<intersection>-148.5 2</intersection>
<intersection>-148 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-148,164.5,-148</points>
<connection>
<GID>326</GID>
<name>set</name></connection>
<connection>
<GID>310</GID>
<name>set</name></connection>
<connection>
<GID>302</GID>
<name>set</name></connection>
<intersection>52.5 5</intersection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-148,111,-147.5</points>
<connection>
<GID>318</GID>
<name>set</name></connection>
<intersection>-148 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-28,-149,-28,-148.5</points>
<connection>
<GID>358</GID>
<name>set</name></connection>
<intersection>-148.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-3,-149,-3,-148.5</points>
<connection>
<GID>350</GID>
<name>set</name></connection>
<intersection>-148.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-160,-55.5,-134</points>
<intersection>-160 2</intersection>
<intersection>-134 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-134,-55.5,-134</points>
<connection>
<GID>366</GID>
<name>OUT_2</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-160,53,-160</points>
<connection>
<GID>336</GID>
<name>set</name></connection>
<intersection>-55.5 0</intersection>
<intersection>-27.5 5</intersection>
<intersection>-2.5 4</intersection>
<intersection>53 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-2.5,-160,-2.5,-159.5</points>
<connection>
<GID>352</GID>
<name>set</name></connection>
<intersection>-160 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-27.5,-160,-27.5,-159.5</points>
<connection>
<GID>360</GID>
<name>set</name></connection>
<intersection>-160 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>53,-160,53,-158.5</points>
<connection>
<GID>344</GID>
<name>set</name></connection>
<intersection>-160 2</intersection>
<intersection>-158.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>53,-158.5,165,-158.5</points>
<connection>
<GID>328</GID>
<name>set</name></connection>
<connection>
<GID>312</GID>
<name>set</name></connection>
<connection>
<GID>304</GID>
<name>set</name></connection>
<intersection>53 7</intersection>
<intersection>111.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>111.5,-158.5,111.5,-158</points>
<connection>
<GID>320</GID>
<name>set</name></connection>
<intersection>-158.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-170.5,-54.5,-135</points>
<intersection>-170.5 2</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-135,-54.5,-135</points>
<connection>
<GID>366</GID>
<name>OUT_1</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54.5,-170.5,52.5,-170.5</points>
<connection>
<GID>362</GID>
<name>set</name></connection>
<connection>
<GID>354</GID>
<name>set</name></connection>
<intersection>-54.5 0</intersection>
<intersection>24 4</intersection>
<intersection>52.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,-171,24,-170.5</points>
<connection>
<GID>338</GID>
<name>set</name></connection>
<intersection>-170.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>52.5,-170.5,52.5,-169.5</points>
<connection>
<GID>346</GID>
<name>set</name></connection>
<intersection>-170.5 2</intersection>
<intersection>-169.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-169.5,164.5,-169.5</points>
<connection>
<GID>330</GID>
<name>set</name></connection>
<connection>
<GID>314</GID>
<name>set</name></connection>
<connection>
<GID>306</GID>
<name>set</name></connection>
<intersection>52.5 5</intersection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-169.5,111,-169</points>
<connection>
<GID>322</GID>
<name>set</name></connection>
<intersection>-169.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-181,-53.5,-136</points>
<intersection>-181 2</intersection>
<intersection>-136 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-136,-53.5,-136</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-181,52.5,-181</points>
<connection>
<GID>364</GID>
<name>set</name></connection>
<connection>
<GID>356</GID>
<name>set</name></connection>
<intersection>-53.5 0</intersection>
<intersection>24 6</intersection>
<intersection>52.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>24,-181.5,24,-181</points>
<connection>
<GID>340</GID>
<name>set</name></connection>
<intersection>-181 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>52.5,-181,52.5,-180</points>
<connection>
<GID>348</GID>
<name>set</name></connection>
<intersection>-181 2</intersection>
<intersection>-180 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>52.5,-180,164.5,-180</points>
<connection>
<GID>332</GID>
<name>set</name></connection>
<connection>
<GID>316</GID>
<name>set</name></connection>
<connection>
<GID>308</GID>
<name>set</name></connection>
<intersection>52.5 7</intersection>
<intersection>111 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>111,-180,111,-179.5</points>
<connection>
<GID>324</GID>
<name>set</name></connection>
<intersection>-180 8</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-183,-34,-106.5</points>
<intersection>-183 1</intersection>
<intersection>-172.5 2</intersection>
<intersection>-161.5 3</intersection>
<intersection>-151 4</intersection>
<intersection>-138.5 5</intersection>
<intersection>-128 6</intersection>
<intersection>-117 7</intersection>
<intersection>-106.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-183,-31,-183</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-172.5,-31,-172.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-34,-161.5,-30.5,-161.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-34,-151,-31,-151</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-34,-138.5,-31,-138.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-34,-128,-31,-128</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-34,-117,-30.5,-117</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-34,-106.5,-31,-106.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection>
<intersection>-33.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-33.5,-106.5,-33.5,-91.5</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>-106.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-183,-11.5,-89.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>-183 1</intersection>
<intersection>-172.5 2</intersection>
<intersection>-161.5 3</intersection>
<intersection>-151 4</intersection>
<intersection>-138.5 5</intersection>
<intersection>-128 6</intersection>
<intersection>-117 7</intersection>
<intersection>-106 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-183,-6,-183</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-172.5,-6,-172.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11.5,-161.5,-5.5,-161.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-11.5,-151,-6,-151</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-11.5,-138.5,-6,-138.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-11.5,-128,-6,-128</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-11.5,-117,-5.5,-117</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-11.5,-106,-5.5,-106</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-183.5,14.5,-89.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>-183.5 1</intersection>
<intersection>-173 2</intersection>
<intersection>-162 3</intersection>
<intersection>-152 4</intersection>
<intersection>-137.5 5</intersection>
<intersection>-127 6</intersection>
<intersection>-116 7</intersection>
<intersection>-105.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-183.5,21,-183.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-173,21,-173</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-162,21.5,-162</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-152,21,-152</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-137.5,20.5,-137.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>14.5,-127,20.5,-127</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>14.5,-116,21,-116</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>14.5,-105.5,20.5,-105.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-182.5,40.5,-104.5</points>
<intersection>-182.5 1</intersection>
<intersection>-172 2</intersection>
<intersection>-161 3</intersection>
<intersection>-150.5 4</intersection>
<intersection>-136.5 5</intersection>
<intersection>-126 6</intersection>
<intersection>-115 7</intersection>
<intersection>-104.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-182.5,49.5,-182.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-172,49.5,-172</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40.5,-161,50,-161</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40.5,-150.5,49.5,-150.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>40.5,-136.5,49,-136.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-126,49.5,-126</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-115,50,-115</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>40,-104.5,49.5,-104.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>40 9</intersection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>40,-104.5,40,-91</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-104.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-182,71,-90.5</points>
<intersection>-182 1</intersection>
<intersection>-171.5 2</intersection>
<intersection>-160.5 3</intersection>
<intersection>-150 4</intersection>
<intersection>-135.5 5</intersection>
<intersection>-125 6</intersection>
<intersection>-114 7</intersection>
<intersection>-103.5 8</intersection>
<intersection>-90.5 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-182,79.5,-182</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-171.5,79.5,-171.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71,-160.5,80.5,-160.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>71,-150,80,-150</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>71,-135.5,81,-135.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>71,-125,81,-125</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>71,-114,81.5,-114</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>71,-103.5,81,-103.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>70.5,-90.5,71,-90.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-181.5,101,-103</points>
<intersection>-181.5 1</intersection>
<intersection>-171 2</intersection>
<intersection>-160 3</intersection>
<intersection>-149.5 4</intersection>
<intersection>-135 5</intersection>
<intersection>-124.5 6</intersection>
<intersection>-113.5 7</intersection>
<intersection>-103 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-181.5,108,-181.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-171,108,-171</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-160,108.5,-160</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101,-149.5,108,-149.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101,-135,108,-135</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>101,-124.5,108,-124.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>101,-113.5,108.5,-113.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>101,-103,108,-103</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection>
<intersection>101.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>101.5,-103,101.5,-94</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>-103 8</intersection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-182,127.5,-92</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-182 1</intersection>
<intersection>-171.5 2</intersection>
<intersection>-160.5 3</intersection>
<intersection>-150 4</intersection>
<intersection>-134.5 5</intersection>
<intersection>-124 6</intersection>
<intersection>-113 9</intersection>
<intersection>-102.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-182,134,-182</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-171.5,134,-171.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127.5,-160.5,134.5,-160.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>127.5,-150,134,-150</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>127.5,-134.5,134.5,-134.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>127.5,-124,134.5,-124</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-102.5,134.5,-102.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>127.5,-113,135,-113</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-182,149.5,-135</points>
<intersection>-182 1</intersection>
<intersection>-135 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-182,161.5,-182</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection>
<intersection>149.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>148.5,-182,148.5,-114</points>
<intersection>-182 1</intersection>
<intersection>-171.5 4</intersection>
<intersection>-160.5 6</intersection>
<intersection>-150 8</intersection>
<intersection>-135 9</intersection>
<intersection>-125 11</intersection>
<intersection>-114 13</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>148.5,-171.5,161.5,-171.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>148.5,-160.5,162,-160.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>148.5,-150,161.5,-150</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>148.5,-135,162.5,-135</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>148.5,-125,163,-125</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>148.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>148,-114,162.5,-114</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>148 14</intersection>
<intersection>148.5 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>148,-114,148,-93.5</points>
<intersection>-114 13</intersection>
<intersection>-103.5 15</intersection>
<intersection>-93.5 16</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>148,-103.5,162.5,-103.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>148 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>146.5,-93.5,148,-93.5</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>148 14</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-72.5,-52,-72.5</points>
<connection>
<GID>376</GID>
<name>CLK</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52.5,-66,-49.5,-66</points>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-134,-69,-132.5</points>
<intersection>-134 1</intersection>
<intersection>-132.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-134,-68,-134</points>
<connection>
<GID>366</GID>
<name>IN_2</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,-132.5,-69,-132.5</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-139.5,-69.5,-136</points>
<intersection>-139.5 2</intersection>
<intersection>-136 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-136,-68,-136</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,-139.5,-69.5,-139.5</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-74,-135,-68,-135</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-195,-22,-112.5</points>
<intersection>-195 4</intersection>
<intersection>-189 11</intersection>
<intersection>-183 12</intersection>
<intersection>-178.5 10</intersection>
<intersection>-167.5 9</intersection>
<intersection>-157 8</intersection>
<intersection>-144.5 7</intersection>
<intersection>-134 6</intersection>
<intersection>-123 5</intersection>
<intersection>-112.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-28,-112.5,-22,-112.5</points>
<connection>
<GID>153</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-24.5,-195,-22,-195</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-27.5,-123,-22,-123</points>
<connection>
<GID>155</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-28,-134,-22,-134</points>
<connection>
<GID>157</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-28,-144.5,-22,-144.5</points>
<connection>
<GID>159</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-28,-157,-22,-157</points>
<connection>
<GID>358</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-27.5,-167.5,-22,-167.5</points>
<connection>
<GID>360</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-28,-178.5,-22,-178.5</points>
<connection>
<GID>362</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-28,-189,-22,-189</points>
<connection>
<GID>364</GID>
<name>clear</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-25,-183,-19.5,-183</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-195,5,-112</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>-189 10</intersection>
<intersection>-178.5 9</intersection>
<intersection>-167.5 8</intersection>
<intersection>-157 7</intersection>
<intersection>-144.5 6</intersection>
<intersection>-134 5</intersection>
<intersection>-123 4</intersection>
<intersection>-112 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2.5,-112,5,-112</points>
<connection>
<GID>161</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-2.5,-123,5,-123</points>
<connection>
<GID>167</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-3,-134,5,-134</points>
<connection>
<GID>170</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-3,-144.5,5,-144.5</points>
<connection>
<GID>176</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-3,-157,5,-157</points>
<connection>
<GID>350</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-2.5,-167.5,5,-167.5</points>
<connection>
<GID>352</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-3,-178.5,5,-178.5</points>
<connection>
<GID>354</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-3,-189,5,-189</points>
<connection>
<GID>356</GID>
<name>clear</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-192.5,31.5,-111.5</points>
<intersection>-192.5 7</intersection>
<intersection>-189.5 4</intersection>
<intersection>-179 5</intersection>
<intersection>-168 6</intersection>
<intersection>-158 8</intersection>
<intersection>-143.5 9</intersection>
<intersection>-133 10</intersection>
<intersection>-122 11</intersection>
<intersection>-111.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-111.5,31.5,-111.5</points>
<connection>
<GID>178</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>24,-189.5,31.5,-189.5</points>
<connection>
<GID>340</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24,-179,31.5,-179</points>
<connection>
<GID>338</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24.5,-168,31.5,-168</points>
<connection>
<GID>336</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>28.5,-192.5,31.5,-192.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>24,-158,31.5,-158</points>
<connection>
<GID>334</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>23.5,-143.5,31.5,-143.5</points>
<connection>
<GID>186</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>23.5,-133,31.5,-133</points>
<connection>
<GID>183</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>24,-122,31.5,-122</points>
<connection>
<GID>180</GID>
<name>clear</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-193,60,-110.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-188.5 4</intersection>
<intersection>-178 5</intersection>
<intersection>-167 6</intersection>
<intersection>-156.5 7</intersection>
<intersection>-142.5 8</intersection>
<intersection>-132 9</intersection>
<intersection>-121 10</intersection>
<intersection>-110.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52.5,-110.5,60,-110.5</points>
<connection>
<GID>211</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-188.5,60,-188.5</points>
<connection>
<GID>348</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>52.5,-178,60,-178</points>
<connection>
<GID>346</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>53,-167,60,-167</points>
<connection>
<GID>344</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>52.5,-156.5,60,-156.5</points>
<connection>
<GID>342</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>52,-142.5,60,-142.5</points>
<connection>
<GID>247</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>52.5,-132,60,-132</points>
<connection>
<GID>219</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>53,-121,60,-121</points>
<connection>
<GID>217</GID>
<name>clear</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-150,92,-109.5</points>
<intersection>-150 2</intersection>
<intersection>-141.5 7</intersection>
<intersection>-131 6</intersection>
<intersection>-120 5</intersection>
<intersection>-109.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91.5,-191,91.5,-150</points>
<intersection>-191 4</intersection>
<intersection>-177.5 10</intersection>
<intersection>-166.5 9</intersection>
<intersection>-156 8</intersection>
<intersection>-150 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-150,92,-150</points>
<intersection>91.5 1</intersection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>84,-109.5,92,-109.5</points>
<connection>
<GID>254</GID>
<name>clear</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-191,91.5,-191</points>
<intersection>82.5 12</intersection>
<intersection>87.5 13</intersection>
<intersection>91.5 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>84.5,-120,92,-120</points>
<connection>
<GID>261</GID>
<name>clear</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>84,-131,92,-131</points>
<connection>
<GID>265</GID>
<name>clear</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>84,-141.5,92,-141.5</points>
<connection>
<GID>269</GID>
<name>clear</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>83,-156,91.5,-156</points>
<connection>
<GID>326</GID>
<name>clear</name></connection>
<intersection>91.5 1</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>83.5,-166.5,91.5,-166.5</points>
<connection>
<GID>328</GID>
<name>clear</name></connection>
<intersection>91.5 1</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>82.5,-177.5,91.5,-177.5</points>
<connection>
<GID>330</GID>
<name>clear</name></connection>
<intersection>91.5 1</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>82.5,-191,82.5,-188</points>
<connection>
<GID>332</GID>
<name>clear</name></connection>
<intersection>-191 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>87.5,-193,87.5,-191</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-191 4</intersection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-192,119.5,-109</points>
<intersection>-192 4</intersection>
<intersection>-177 10</intersection>
<intersection>-166 9</intersection>
<intersection>-155.5 8</intersection>
<intersection>-141 7</intersection>
<intersection>-130.5 6</intersection>
<intersection>-119.5 5</intersection>
<intersection>-109 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>111,-109,119.5,-109</points>
<connection>
<GID>273</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-192,119.5,-192</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>111 11</intersection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>111.5,-119.5,119.5,-119.5</points>
<connection>
<GID>277</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>111,-130.5,119.5,-130.5</points>
<connection>
<GID>281</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>111,-141,119.5,-141</points>
<connection>
<GID>284</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>111,-155.5,119.5,-155.5</points>
<connection>
<GID>318</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>111.5,-166,119.5,-166</points>
<connection>
<GID>320</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>111,-177,119.5,-177</points>
<connection>
<GID>322</GID>
<name>clear</name></connection>
<intersection>119.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>111,-192,111,-187.5</points>
<connection>
<GID>324</GID>
<name>clear</name></connection>
<intersection>-192 4</intersection></vsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-192.5,146,-108.5</points>
<intersection>-192.5 4</intersection>
<intersection>-177.5 10</intersection>
<intersection>-166.5 9</intersection>
<intersection>-156 8</intersection>
<intersection>-140.5 7</intersection>
<intersection>-130 6</intersection>
<intersection>-119 5</intersection>
<intersection>-108.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>137.5,-108.5,146,-108.5</points>
<connection>
<GID>286</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>137,-192.5,146,-192.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>137 11</intersection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>138,-119,146,-119</points>
<connection>
<GID>288</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>137.5,-130,146,-130</points>
<connection>
<GID>290</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>137.5,-140.5,146,-140.5</points>
<connection>
<GID>292</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>137,-156,146,-156</points>
<connection>
<GID>310</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>137.5,-166.5,146,-166.5</points>
<connection>
<GID>312</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>137,-177.5,146,-177.5</points>
<connection>
<GID>314</GID>
<name>clear</name></connection>
<intersection>146 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>137,-192.5,137,-188</points>
<connection>
<GID>316</GID>
<name>clear</name></connection>
<intersection>-192.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-193,175.5,-109.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-177.5 9</intersection>
<intersection>-166.5 8</intersection>
<intersection>-156 7</intersection>
<intersection>-141 6</intersection>
<intersection>-131 5</intersection>
<intersection>-120 4</intersection>
<intersection>-109.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>165.5,-109.5,175.5,-109.5</points>
<connection>
<GID>294</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>165.5,-120,175.5,-120</points>
<connection>
<GID>296</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>166,-131,175.5,-131</points>
<connection>
<GID>298</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>165.5,-141,175.5,-141</points>
<connection>
<GID>300</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>164.5,-156,175.5,-156</points>
<connection>
<GID>302</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>165,-166.5,175.5,-166.5</points>
<connection>
<GID>304</GID>
<name>clear</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>164.5,-177.5,175.5,-177.5</points>
<connection>
<GID>306</GID>
<name>clear</name></connection>
<intersection>174 12</intersection>
<intersection>175.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>174,-188,174,-177.5</points>
<intersection>-188 13</intersection>
<intersection>-177.5 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>164.5,-188,174,-188</points>
<connection>
<GID>308</GID>
<name>clear</name></connection>
<intersection>174 12</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-106.5,-24,-106</points>
<intersection>-106.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-106.5,-24,-106.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24,-106,-23,-106</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-117.5,-22.5,-117</points>
<intersection>-117.5 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-117,-22.5,-117</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,-117.5,-20,-117.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-128,-21,-128</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-139.5,-23,-138.5</points>
<intersection>-139.5 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-138.5,-23,-138.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-139.5,-21,-139.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-151,-21,-151</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-162.5,-23,-161.5</points>
<intersection>-162.5 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-161.5,-23,-161.5</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-162.5,-21.5,-162.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-173,-23,-172.5</points>
<intersection>-173 2</intersection>
<intersection>-172.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-172.5,-23,-172.5</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,-173,-21,-173</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-106,3.5,-106</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<connection>
<GID>399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-117,2,-117</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-128.5,0.5,-128</points>
<intersection>-128.5 1</intersection>
<intersection>-128 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-128.5,1.5,-128.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-128,0.5,-128</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-138.5,2.5,-138.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-151,1,-150.5</points>
<intersection>-151 1</intersection>
<intersection>-150.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-151,1,-151</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-150.5,2,-150.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-161.5,2,-161.5</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<connection>
<GID>404</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-173,0.5,-172.5</points>
<intersection>-173 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-173,1.5,-173</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-172.5,0.5,-172.5</points>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-183.5,0.5,-183</points>
<intersection>-183.5 2</intersection>
<intersection>-183 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-183,0.5,-183</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0.5,-183.5,1.5,-183.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-105.5,27.5,-104.5</points>
<intersection>-105.5 1</intersection>
<intersection>-104.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-105.5,27.5,-105.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-104.5,29,-104.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-116,28.5,-116</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-127,27.5,-126</points>
<intersection>-127 1</intersection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-127,27.5,-127</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-126,29,-126</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-137.5,27.5,-137</points>
<intersection>-137.5 1</intersection>
<intersection>-137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-137.5,27.5,-137.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-137,29,-137</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-152,28,-151.5</points>
<intersection>-152 2</intersection>
<intersection>-151.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-151.5,29,-151.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-152,28,-152</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-162,29.5,-162</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<connection>
<GID>412</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-173,28,-172.5</points>
<intersection>-173 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-173,28,-173</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-172.5,29.5,-172.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-183.5,30,-183.5</points>
<connection>
<GID>340</GID>
<name>OUT_0</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-105,57,-104.5</points>
<intersection>-105 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-104.5,57,-104.5</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-105,59,-105</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-115,58,-115</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-126,58.5,-126</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<connection>
<GID>417</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-136.5,58,-136.5</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<connection>
<GID>418</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-151,56.5,-150.5</points>
<intersection>-151 2</intersection>
<intersection>-150.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-150.5,56.5,-150.5</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-151,57.5,-151</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-161,57,-160.5</points>
<intersection>-161 1</intersection>
<intersection>-160.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-161,57,-161</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-160.5,58,-160.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-172,56.5,-171.5</points>
<intersection>-172 1</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-172,56.5,-172</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-171.5,58,-171.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-182.5,56.5,-181.5</points>
<intersection>-182.5 1</intersection>
<intersection>-181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-182.5,56.5,-182.5</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-181.5,57.5,-181.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-105,88,-103.5</points>
<intersection>-105 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-103.5,88,-103.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88,-105,89,-105</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-114,90,-114</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<connection>
<GID>424</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-125,88.5,-124.5</points>
<intersection>-125 1</intersection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-125,88.5,-125</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-124.5,90.5,-124.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-135.5,89.5,-135.5</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<connection>
<GID>426</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-150,87.5,-149.5</points>
<intersection>-150 1</intersection>
<intersection>-149.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-150,87.5,-150</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-149.5,89.5,-149.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-160.5,87.5,-160</points>
<intersection>-160.5 1</intersection>
<intersection>-160 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-160.5,87.5,-160.5</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-160,88.5,-160</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-171.5,87,-171</points>
<intersection>-171.5 1</intersection>
<intersection>-171 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-171.5,87,-171.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-171,89,-171</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-182,87,-181.5</points>
<intersection>-182 1</intersection>
<intersection>-181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-182,87,-182</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-181.5,88.5,-181.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-103.5,115,-103</points>
<intersection>-103.5 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-103,115,-103</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-103.5,116,-103.5</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,-113.5,116.5,-113.5</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<connection>
<GID>432</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-125,114.5,-124.5</points>
<intersection>-125 1</intersection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-125,115,-125</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-124.5,114.5,-124.5</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-137,115,-135</points>
<intersection>-137 2</intersection>
<intersection>-135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-135,115,-135</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-137,116.5,-137</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-149.5,115,-149</points>
<intersection>-149.5 1</intersection>
<intersection>-149 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-149.5,115,-149.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-149,116.5,-149</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,-160,115.5,-160</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<connection>
<GID>436</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-171.5,115,-171</points>
<intersection>-171.5 1</intersection>
<intersection>-171 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-171.5,116,-171.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-171,115,-171</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-181.5,115,-181</points>
<intersection>-181.5 1</intersection>
<intersection>-181 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-181.5,115,-181.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-181,116,-181</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-104,141,-102.5</points>
<intersection>-104 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-102.5,141,-102.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-104,141.5,-104</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-113.5,142,-113</points>
<intersection>-113.5 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-113.5,143,-113.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-113,142,-113</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-124.5,141.5,-124</points>
<intersection>-124.5 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-124.5,142.5,-124.5</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-124,141.5,-124</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-135,141.5,-134.5</points>
<intersection>-135 1</intersection>
<intersection>-134.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-135,142.5,-135</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-134.5,141.5,-134.5</points>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-150.5,141,-150</points>
<intersection>-150.5 1</intersection>
<intersection>-150 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-150.5,142,-150.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-150,141,-150</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-161,141,-160.5</points>
<intersection>-161 1</intersection>
<intersection>-160.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-161,142,-161</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-160.5,141,-160.5</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-172.5,140.5,-171.5</points>
<intersection>-172.5 1</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-172.5,141.5,-172.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-171.5,140.5,-171.5</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-184,141,-182</points>
<intersection>-184 2</intersection>
<intersection>-182 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-182,141,-182</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-184,142,-184</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-103.5,170.5,-103</points>
<intersection>-103.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-103.5,170.5,-103.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-103,173,-103</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168.5,-114,172.5,-114</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169,-125,171.5,-125</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168.5,-135,172,-135</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-150,172,-150</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-161,170,-160.5</points>
<intersection>-161 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-160.5,170,-160.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-161,172,-161</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-171.5,171.5,-171.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-182,171.5,-182</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-71.5,78.5,-66.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>444</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-71.5,84.5,-66.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-72,90,-66.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-71.5,95.5,-66.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-71.5,101,-66.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>448</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-72,106.5,-68</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>449</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-72,112,-66.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-71.5,117.5,-66.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<connection>
<GID>451</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158.5,-66.5,169.5,-66.5</points>
<connection>
<GID>181</GID>
<name>IN_7</name></connection>
<intersection>158.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158.5,-66.5,158.5,-66</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>-66.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-68.5,161,-67.5</points>
<intersection>-68.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-67.5,169.5,-67.5</points>
<connection>
<GID>181</GID>
<name>IN_6</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-68.5,161,-68.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-71,160,-68.5</points>
<intersection>-71 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-68.5,169.5,-68.5</points>
<connection>
<GID>181</GID>
<name>IN_5</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>158,-71,160,-71</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-75,160.5,-69.5</points>
<intersection>-75 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-69.5,169.5,-69.5</points>
<connection>
<GID>181</GID>
<name>IN_4</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,-75,160.5,-75</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-79,161,-70.5</points>
<intersection>-79 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-70.5,169.5,-70.5</points>
<connection>
<GID>181</GID>
<name>IN_3</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-79,161,-79</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-82,163,-71.5</points>
<intersection>-82 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-71.5,169.5,-71.5</points>
<connection>
<GID>181</GID>
<name>IN_2</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-82,163,-82</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-85,164.5,-72.5</points>
<intersection>-85 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-72.5,169.5,-72.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>164.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>164.5,-85,165,-85</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-80,168.5,-73.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-73.5,169.5,-73.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-202,113,-202</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>113 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>113,-204,113,-202</points>
<connection>
<GID>471</GID>
<name>IN_7</name></connection>
<intersection>-202 1</intersection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-205,113,-205</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>113 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>113,-205,113,-205</points>
<connection>
<GID>471</GID>
<name>IN_6</name></connection>
<intersection>-205 1</intersection></vsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-205.5,113,-205.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113,-206,113,-205.5</points>
<connection>
<GID>471</GID>
<name>IN_5</name></connection>
<intersection>-205.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-207.5,110.5,-207</points>
<intersection>-207.5 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-207,113,-207</points>
<connection>
<GID>471</GID>
<name>IN_4</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-207.5,110.5,-207.5</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100,-208.5,113,-208.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>113 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>113,-208.5,113,-208</points>
<connection>
<GID>471</GID>
<name>IN_3</name></connection>
<intersection>-208.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-210,110.5,-209</points>
<intersection>-210 2</intersection>
<intersection>-209 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-209,113,-209</points>
<connection>
<GID>471</GID>
<name>IN_2</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-210,110.5,-210</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-213,111,-210</points>
<intersection>-213 2</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-210,113,-210</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-213,111,-213</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-216,113,-211</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>-216 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110.5,-216,113,-216</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,-222,113.5,-222</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113.5,-224,113.5,-222</points>
<connection>
<GID>482</GID>
<name>IN_7</name></connection>
<intersection>-222 1</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-224.5,113.5,-224.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>113.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>113.5,-225,113.5,-224.5</points>
<connection>
<GID>482</GID>
<name>IN_6</name></connection>
<intersection>-224.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102,-226,113.5,-226</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>113.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113.5,-226,113.5,-226</points>
<connection>
<GID>482</GID>
<name>IN_5</name></connection>
<intersection>-226 1</intersection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-227.5,111,-227</points>
<intersection>-227.5 2</intersection>
<intersection>-227 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-227,113.5,-227</points>
<connection>
<GID>482</GID>
<name>IN_4</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-227.5,111,-227.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98.5,-229,113.5,-229</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113.5,-229,113.5,-228</points>
<connection>
<GID>482</GID>
<name>IN_3</name></connection>
<intersection>-229 1</intersection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-230,111,-229</points>
<intersection>-230 2</intersection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-229,113.5,-229</points>
<connection>
<GID>482</GID>
<name>IN_2</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-230,111,-230</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-233,111.5,-230</points>
<intersection>-233 2</intersection>
<intersection>-230 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-230,113.5,-230</points>
<connection>
<GID>482</GID>
<name>IN_1</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-233,111.5,-233</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-236,113.5,-231</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-236 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-236,114,-236</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113,-242,114,-242</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>114 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114,-242,114,-242</points>
<connection>
<GID>491</GID>
<name>IN_7</name></connection>
<intersection>-242 1</intersection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-243.5,114,-243.5</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>114 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114,-243.5,114,-243</points>
<connection>
<GID>491</GID>
<name>IN_6</name></connection>
<intersection>-243.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,-240.5,114,-240.5</points>
<intersection>97.5 5</intersection>
<intersection>114 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114,-244,114,-240.5</points>
<connection>
<GID>491</GID>
<name>IN_5</name></connection>
<intersection>-240.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>97.5,-243,97.5,-240.5</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-240.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-245.5,111.5,-245</points>
<intersection>-245.5 2</intersection>
<intersection>-245 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-245,114,-245</points>
<connection>
<GID>491</GID>
<name>IN_4</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-245.5,111.5,-245.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,-246.5,114,-246.5</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>114 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114,-246.5,114,-246</points>
<connection>
<GID>491</GID>
<name>IN_3</name></connection>
<intersection>-246.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-248.5,111.5,-247</points>
<intersection>-248.5 2</intersection>
<intersection>-247 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-247,114,-247</points>
<connection>
<GID>491</GID>
<name>IN_2</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-248.5,111.5,-248.5</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-251,112,-248</points>
<intersection>-251 2</intersection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-248,114,-248</points>
<connection>
<GID>491</GID>
<name>IN_1</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-251,112,-251</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-254,114,-249</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-254 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-254,114.5,-254</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113,-258.5,114,-258.5</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>114 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114,-258.5,114,-258.5</points>
<connection>
<GID>500</GID>
<name>IN_7</name></connection>
<intersection>-258.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-259.5,114,-259.5</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>114 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114,-259.5,114,-259.5</points>
<connection>
<GID>500</GID>
<name>IN_6</name></connection>
<intersection>-259.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-260.5,114,-260.5</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>114 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>114,-260.5,114,-260.5</points>
<connection>
<GID>500</GID>
<name>IN_5</name></connection>
<intersection>-260.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-262,111.5,-261.5</points>
<intersection>-262 2</intersection>
<intersection>-261.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-261.5,114,-261.5</points>
<connection>
<GID>500</GID>
<name>IN_4</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-262,111.5,-262</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101.5,-263.5,114,-263.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>114 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114,-263.5,114,-262.5</points>
<connection>
<GID>500</GID>
<name>IN_3</name></connection>
<intersection>-263.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-264.5,111.5,-263.5</points>
<intersection>-264.5 2</intersection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-263.5,114,-263.5</points>
<connection>
<GID>500</GID>
<name>IN_2</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-264.5,111.5,-264.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-267.5,112,-264.5</points>
<intersection>-267.5 2</intersection>
<intersection>-264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-264.5,114,-264.5</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-267.5,112,-267.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-270.5,114,-265.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-270.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-270.5,114.5,-270.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,-275.5,114.5,-275.5</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>114.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-277,114.5,-275.5</points>
<connection>
<GID>509</GID>
<name>IN_7</name></connection>
<intersection>-275.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,-278,114.5,-278</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-278,114.5,-278</points>
<connection>
<GID>509</GID>
<name>IN_6</name></connection>
<intersection>-278 1</intersection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-279,114.5,-279</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-279,114.5,-279</points>
<connection>
<GID>509</GID>
<name>IN_5</name></connection>
<intersection>-279 1</intersection></vsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-280.5,112,-280</points>
<intersection>-280.5 2</intersection>
<intersection>-280 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-280,114.5,-280</points>
<connection>
<GID>509</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-280.5,112,-280.5</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102.5,-281,114.5,-281</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>114.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>114.5,-281,114.5,-281</points>
<connection>
<GID>509</GID>
<name>IN_3</name></connection>
<intersection>-281 1</intersection></vsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-283,112,-282</points>
<intersection>-283 2</intersection>
<intersection>-282 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-282,114.5,-282</points>
<connection>
<GID>509</GID>
<name>IN_2</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-283,112,-283</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-286,112.5,-283</points>
<intersection>-286 2</intersection>
<intersection>-283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-283,114.5,-283</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-286,112.5,-286</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-289,114.5,-284</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-289,115,-289</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-296.5,114.5,-296.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-296.5,114.5,-296.5</points>
<connection>
<GID>518</GID>
<name>IN_7</name></connection>
<intersection>-296.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,-297.5,114.5,-297.5</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-297.5,114.5,-297.5</points>
<connection>
<GID>518</GID>
<name>IN_6</name></connection>
<intersection>-297.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-298,114.5,-298</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>114.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-298.5,114.5,-298</points>
<connection>
<GID>518</GID>
<name>IN_5</name></connection>
<intersection>-298 1</intersection></vsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-300,112,-299.5</points>
<intersection>-300 2</intersection>
<intersection>-299.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-299.5,114.5,-299.5</points>
<connection>
<GID>518</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-300,112,-300</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-301,114.5,-301</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>114.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-301,114.5,-300.5</points>
<connection>
<GID>518</GID>
<name>IN_3</name></connection>
<intersection>-301 1</intersection></vsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-302.5,112,-301.5</points>
<intersection>-302.5 2</intersection>
<intersection>-301.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-301.5,114.5,-301.5</points>
<connection>
<GID>518</GID>
<name>IN_2</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-302.5,112,-302.5</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-305.5,112.5,-302.5</points>
<intersection>-305.5 2</intersection>
<intersection>-302.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-302.5,114.5,-302.5</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-305.5,112.5,-305.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-308.5,114.5,-303.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>-308.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-308.5,115,-308.5</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-315.5,114.5,-315.5</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>114.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-316.5,114.5,-315.5</points>
<connection>
<GID>527</GID>
<name>IN_7</name></connection>
<intersection>-315.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,-317.5,114.5,-317.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-317.5,114.5,-317.5</points>
<connection>
<GID>527</GID>
<name>IN_6</name></connection>
<intersection>-317.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-318.5,114.5,-318.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-318.5,114.5,-318.5</points>
<connection>
<GID>527</GID>
<name>IN_5</name></connection>
<intersection>-318.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-320,112,-319.5</points>
<intersection>-320 2</intersection>
<intersection>-319.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-319.5,114.5,-319.5</points>
<connection>
<GID>527</GID>
<name>IN_4</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-320,112,-320</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98.5,-320.5,114.5,-320.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>114.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>114.5,-320.5,114.5,-320.5</points>
<connection>
<GID>527</GID>
<name>IN_3</name></connection>
<intersection>-320.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-322.5,112,-321.5</points>
<intersection>-322.5 2</intersection>
<intersection>-321.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-321.5,114.5,-321.5</points>
<connection>
<GID>527</GID>
<name>IN_2</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-322.5,112,-322.5</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-325.5,112.5,-322.5</points>
<intersection>-325.5 2</intersection>
<intersection>-322.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-322.5,114.5,-322.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-325.5,112.5,-325.5</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-328.5,114.5,-323.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-328.5,115,-328.5</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,-335,115.5,-335</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>115.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>115.5,-335,115.5,-335</points>
<connection>
<GID>536</GID>
<name>IN_7</name></connection>
<intersection>-335 1</intersection></vsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105.5,-334.5,115.5,-334.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>115.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>115.5,-336,115.5,-334.5</points>
<connection>
<GID>536</GID>
<name>IN_6</name></connection>
<intersection>-334.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-337,115.5,-337</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>115.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>115.5,-337,115.5,-337</points>
<connection>
<GID>536</GID>
<name>IN_5</name></connection>
<intersection>-337 1</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-338.5,113,-338</points>
<intersection>-338.5 2</intersection>
<intersection>-338 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-338,115.5,-338</points>
<connection>
<GID>536</GID>
<name>IN_4</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-338.5,113,-338.5</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-339.5,115.5,-339.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>115.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>115.5,-339.5,115.5,-339</points>
<connection>
<GID>536</GID>
<name>IN_3</name></connection>
<intersection>-339.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-341,113,-340</points>
<intersection>-341 2</intersection>
<intersection>-340 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-340,115.5,-340</points>
<connection>
<GID>536</GID>
<name>IN_2</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-341,113,-341</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-344,113.5,-341</points>
<intersection>-344 2</intersection>
<intersection>-341 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-341,115.5,-341</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-344,113.5,-344</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-347,115.5,-342</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>-347 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-347,116,-347</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 1>
<page 2>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 2>
<page 3>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 3>
<page 4>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 4>
<page 5>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 5>
<page 6>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 6>
<page 7>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 7>
<page 8>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 8>
<page 9>
<PageViewport>-1e+010,105.438,-1e+010,-491.562</PageViewport></page 9></circuit>